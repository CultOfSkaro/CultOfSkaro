-------------------------------------------------------------------------------
-- plb_bram_if_cntlr_1_bram_elaborate.vhd
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

entity plb_bram_if_cntlr_1_bram_elaborate is
  generic (
    C_MEMSIZE : integer;
    C_PORT_DWIDTH : integer;
    C_PORT_AWIDTH : integer;
    C_NUM_WE : integer;
    C_FAMILY : string
    );
  port (
    BRAM_Rst_A : in std_logic;
    BRAM_Clk_A : in std_logic;
    BRAM_EN_A : in std_logic;
    BRAM_WEN_A : in std_logic_vector(0 to C_NUM_WE-1);
    BRAM_Addr_A : in std_logic_vector(0 to C_PORT_AWIDTH-1);
    BRAM_Din_A : out std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Dout_A : in std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Rst_B : in std_logic;
    BRAM_Clk_B : in std_logic;
    BRAM_EN_B : in std_logic;
    BRAM_WEN_B : in std_logic_vector(0 to C_NUM_WE-1);
    BRAM_Addr_B : in std_logic_vector(0 to C_PORT_AWIDTH-1);
    BRAM_Din_B : out std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Dout_B : in std_logic_vector(0 to C_PORT_DWIDTH-1)
  );

  attribute keep_hierarchy : STRING;
  attribute keep_hierarchy of plb_bram_if_cntlr_1_bram_elaborate : entity is "yes";

end plb_bram_if_cntlr_1_bram_elaborate;

architecture STRUCTURE of plb_bram_if_cntlr_1_bram_elaborate is

  component RAMB16 is
    generic (
      WRITE_MODE_A : string;
      WRITE_MODE_B : string;
      INIT_FILE : string;
      READ_WIDTH_A : integer;
      READ_WIDTH_B : integer;
      WRITE_WIDTH_A : integer;
      WRITE_WIDTH_B : integer;
      RAM_EXTENSION_A : string;
      RAM_EXTENSION_B : string
    );
    port (
      ADDRA : in std_logic_vector(14 downto 0);
      CASCADEINA : in std_logic;
      CASCADEOUTA : out std_logic;
      CLKA : in std_logic;
      DIA : in std_logic_vector(31 downto 0);
      DIPA : in std_logic_vector(3 downto 0);
      DOA : out std_logic_vector(31 downto 0);
      DOPA : out std_logic_vector(3 downto 0);
      ENA : in std_logic;
      REGCEA : in std_logic;
      SSRA : in std_logic;
      WEA : in std_logic_vector(3 downto 0);
      ADDRB : in std_logic_vector(14 downto 0);
      CASCADEINB : in std_logic;
      CASCADEOUTB : out std_logic;
      CLKB : in std_logic;
      DIB : in std_logic_vector(31 downto 0);
      DIPB : in std_logic_vector(3 downto 0);
      DOB : out std_logic_vector(31 downto 0);
      DOPB : out std_logic_vector(3 downto 0);
      ENB : in std_logic;
      REGCEB : in std_logic;
      SSRB : in std_logic;
      WEB : in std_logic_vector(3 downto 0)
    );
  end component;

  attribute BMM_INFO : STRING;

  attribute BMM_INFO of ramb16_0: label is " ";
  attribute BMM_INFO of ramb16_1: label is " ";
  attribute BMM_INFO of ramb16_2: label is " ";
  attribute BMM_INFO of ramb16_3: label is " ";
  attribute BMM_INFO of ramb16_4: label is " ";
  attribute BMM_INFO of ramb16_5: label is " ";
  attribute BMM_INFO of ramb16_6: label is " ";
  attribute BMM_INFO of ramb16_7: label is " ";
  attribute BMM_INFO of ramb16_8: label is " ";
  attribute BMM_INFO of ramb16_9: label is " ";
  attribute BMM_INFO of ramb16_10: label is " ";
  attribute BMM_INFO of ramb16_11: label is " ";
  attribute BMM_INFO of ramb16_12: label is " ";
  attribute BMM_INFO of ramb16_13: label is " ";
  attribute BMM_INFO of ramb16_14: label is " ";
  attribute BMM_INFO of ramb16_15: label is " ";
  attribute BMM_INFO of ramb16_16: label is " ";
  attribute BMM_INFO of ramb16_17: label is " ";
  attribute BMM_INFO of ramb16_18: label is " ";
  attribute BMM_INFO of ramb16_19: label is " ";
  attribute BMM_INFO of ramb16_20: label is " ";
  attribute BMM_INFO of ramb16_21: label is " ";
  attribute BMM_INFO of ramb16_22: label is " ";
  attribute BMM_INFO of ramb16_23: label is " ";
  attribute BMM_INFO of ramb16_24: label is " ";
  attribute BMM_INFO of ramb16_25: label is " ";
  attribute BMM_INFO of ramb16_26: label is " ";
  attribute BMM_INFO of ramb16_27: label is " ";
  attribute BMM_INFO of ramb16_28: label is " ";
  attribute BMM_INFO of ramb16_29: label is " ";
  attribute BMM_INFO of ramb16_30: label is " ";
  attribute BMM_INFO of ramb16_31: label is " ";
  attribute BMM_INFO of ramb16_32: label is " ";
  attribute BMM_INFO of ramb16_33: label is " ";
  attribute BMM_INFO of ramb16_34: label is " ";
  attribute BMM_INFO of ramb16_35: label is " ";
  attribute BMM_INFO of ramb16_36: label is " ";
  attribute BMM_INFO of ramb16_37: label is " ";
  attribute BMM_INFO of ramb16_38: label is " ";
  attribute BMM_INFO of ramb16_39: label is " ";
  attribute BMM_INFO of ramb16_40: label is " ";
  attribute BMM_INFO of ramb16_41: label is " ";
  attribute BMM_INFO of ramb16_42: label is " ";
  attribute BMM_INFO of ramb16_43: label is " ";
  attribute BMM_INFO of ramb16_44: label is " ";
  attribute BMM_INFO of ramb16_45: label is " ";
  attribute BMM_INFO of ramb16_46: label is " ";
  attribute BMM_INFO of ramb16_47: label is " ";
  attribute BMM_INFO of ramb16_48: label is " ";
  attribute BMM_INFO of ramb16_49: label is " ";
  attribute BMM_INFO of ramb16_50: label is " ";
  attribute BMM_INFO of ramb16_51: label is " ";
  attribute BMM_INFO of ramb16_52: label is " ";
  attribute BMM_INFO of ramb16_53: label is " ";
  attribute BMM_INFO of ramb16_54: label is " ";
  attribute BMM_INFO of ramb16_55: label is " ";
  attribute BMM_INFO of ramb16_56: label is " ";
  attribute BMM_INFO of ramb16_57: label is " ";
  attribute BMM_INFO of ramb16_58: label is " ";
  attribute BMM_INFO of ramb16_59: label is " ";
  attribute BMM_INFO of ramb16_60: label is " ";
  attribute BMM_INFO of ramb16_61: label is " ";
  attribute BMM_INFO of ramb16_62: label is " ";
  attribute BMM_INFO of ramb16_63: label is " ";
  -- Internal signals

  signal net_gnd0 : std_logic;
  signal net_gnd4 : std_logic_vector(3 downto 0);
  signal pgassign1 : std_logic_vector(0 to 0);
  signal pgassign2 : std_logic_vector(0 to 30);
  signal pgassign3 : std_logic_vector(14 downto 0);
  signal pgassign4 : std_logic_vector(31 downto 0);
  signal pgassign5 : std_logic_vector(31 downto 0);
  signal pgassign6 : std_logic_vector(3 downto 0);
  signal pgassign7 : std_logic_vector(14 downto 0);
  signal pgassign8 : std_logic_vector(31 downto 0);
  signal pgassign9 : std_logic_vector(31 downto 0);
  signal pgassign10 : std_logic_vector(3 downto 0);
  signal pgassign11 : std_logic_vector(14 downto 0);
  signal pgassign12 : std_logic_vector(31 downto 0);
  signal pgassign13 : std_logic_vector(31 downto 0);
  signal pgassign14 : std_logic_vector(3 downto 0);
  signal pgassign15 : std_logic_vector(14 downto 0);
  signal pgassign16 : std_logic_vector(31 downto 0);
  signal pgassign17 : std_logic_vector(31 downto 0);
  signal pgassign18 : std_logic_vector(3 downto 0);
  signal pgassign19 : std_logic_vector(14 downto 0);
  signal pgassign20 : std_logic_vector(31 downto 0);
  signal pgassign21 : std_logic_vector(31 downto 0);
  signal pgassign22 : std_logic_vector(3 downto 0);
  signal pgassign23 : std_logic_vector(14 downto 0);
  signal pgassign24 : std_logic_vector(31 downto 0);
  signal pgassign25 : std_logic_vector(31 downto 0);
  signal pgassign26 : std_logic_vector(3 downto 0);
  signal pgassign27 : std_logic_vector(14 downto 0);
  signal pgassign28 : std_logic_vector(31 downto 0);
  signal pgassign29 : std_logic_vector(31 downto 0);
  signal pgassign30 : std_logic_vector(3 downto 0);
  signal pgassign31 : std_logic_vector(14 downto 0);
  signal pgassign32 : std_logic_vector(31 downto 0);
  signal pgassign33 : std_logic_vector(31 downto 0);
  signal pgassign34 : std_logic_vector(3 downto 0);
  signal pgassign35 : std_logic_vector(14 downto 0);
  signal pgassign36 : std_logic_vector(31 downto 0);
  signal pgassign37 : std_logic_vector(31 downto 0);
  signal pgassign38 : std_logic_vector(3 downto 0);
  signal pgassign39 : std_logic_vector(14 downto 0);
  signal pgassign40 : std_logic_vector(31 downto 0);
  signal pgassign41 : std_logic_vector(31 downto 0);
  signal pgassign42 : std_logic_vector(3 downto 0);
  signal pgassign43 : std_logic_vector(14 downto 0);
  signal pgassign44 : std_logic_vector(31 downto 0);
  signal pgassign45 : std_logic_vector(31 downto 0);
  signal pgassign46 : std_logic_vector(3 downto 0);
  signal pgassign47 : std_logic_vector(14 downto 0);
  signal pgassign48 : std_logic_vector(31 downto 0);
  signal pgassign49 : std_logic_vector(31 downto 0);
  signal pgassign50 : std_logic_vector(3 downto 0);
  signal pgassign51 : std_logic_vector(14 downto 0);
  signal pgassign52 : std_logic_vector(31 downto 0);
  signal pgassign53 : std_logic_vector(31 downto 0);
  signal pgassign54 : std_logic_vector(3 downto 0);
  signal pgassign55 : std_logic_vector(14 downto 0);
  signal pgassign56 : std_logic_vector(31 downto 0);
  signal pgassign57 : std_logic_vector(31 downto 0);
  signal pgassign58 : std_logic_vector(3 downto 0);
  signal pgassign59 : std_logic_vector(14 downto 0);
  signal pgassign60 : std_logic_vector(31 downto 0);
  signal pgassign61 : std_logic_vector(31 downto 0);
  signal pgassign62 : std_logic_vector(3 downto 0);
  signal pgassign63 : std_logic_vector(14 downto 0);
  signal pgassign64 : std_logic_vector(31 downto 0);
  signal pgassign65 : std_logic_vector(31 downto 0);
  signal pgassign66 : std_logic_vector(3 downto 0);
  signal pgassign67 : std_logic_vector(14 downto 0);
  signal pgassign68 : std_logic_vector(31 downto 0);
  signal pgassign69 : std_logic_vector(31 downto 0);
  signal pgassign70 : std_logic_vector(3 downto 0);
  signal pgassign71 : std_logic_vector(14 downto 0);
  signal pgassign72 : std_logic_vector(31 downto 0);
  signal pgassign73 : std_logic_vector(31 downto 0);
  signal pgassign74 : std_logic_vector(3 downto 0);
  signal pgassign75 : std_logic_vector(14 downto 0);
  signal pgassign76 : std_logic_vector(31 downto 0);
  signal pgassign77 : std_logic_vector(31 downto 0);
  signal pgassign78 : std_logic_vector(3 downto 0);
  signal pgassign79 : std_logic_vector(14 downto 0);
  signal pgassign80 : std_logic_vector(31 downto 0);
  signal pgassign81 : std_logic_vector(31 downto 0);
  signal pgassign82 : std_logic_vector(3 downto 0);
  signal pgassign83 : std_logic_vector(14 downto 0);
  signal pgassign84 : std_logic_vector(31 downto 0);
  signal pgassign85 : std_logic_vector(31 downto 0);
  signal pgassign86 : std_logic_vector(3 downto 0);
  signal pgassign87 : std_logic_vector(14 downto 0);
  signal pgassign88 : std_logic_vector(31 downto 0);
  signal pgassign89 : std_logic_vector(31 downto 0);
  signal pgassign90 : std_logic_vector(3 downto 0);
  signal pgassign91 : std_logic_vector(14 downto 0);
  signal pgassign92 : std_logic_vector(31 downto 0);
  signal pgassign93 : std_logic_vector(31 downto 0);
  signal pgassign94 : std_logic_vector(3 downto 0);
  signal pgassign95 : std_logic_vector(14 downto 0);
  signal pgassign96 : std_logic_vector(31 downto 0);
  signal pgassign97 : std_logic_vector(31 downto 0);
  signal pgassign98 : std_logic_vector(3 downto 0);
  signal pgassign99 : std_logic_vector(14 downto 0);
  signal pgassign100 : std_logic_vector(31 downto 0);
  signal pgassign101 : std_logic_vector(31 downto 0);
  signal pgassign102 : std_logic_vector(3 downto 0);
  signal pgassign103 : std_logic_vector(14 downto 0);
  signal pgassign104 : std_logic_vector(31 downto 0);
  signal pgassign105 : std_logic_vector(31 downto 0);
  signal pgassign106 : std_logic_vector(3 downto 0);
  signal pgassign107 : std_logic_vector(14 downto 0);
  signal pgassign108 : std_logic_vector(31 downto 0);
  signal pgassign109 : std_logic_vector(31 downto 0);
  signal pgassign110 : std_logic_vector(3 downto 0);
  signal pgassign111 : std_logic_vector(14 downto 0);
  signal pgassign112 : std_logic_vector(31 downto 0);
  signal pgassign113 : std_logic_vector(31 downto 0);
  signal pgassign114 : std_logic_vector(3 downto 0);
  signal pgassign115 : std_logic_vector(14 downto 0);
  signal pgassign116 : std_logic_vector(31 downto 0);
  signal pgassign117 : std_logic_vector(31 downto 0);
  signal pgassign118 : std_logic_vector(3 downto 0);
  signal pgassign119 : std_logic_vector(14 downto 0);
  signal pgassign120 : std_logic_vector(31 downto 0);
  signal pgassign121 : std_logic_vector(31 downto 0);
  signal pgassign122 : std_logic_vector(3 downto 0);
  signal pgassign123 : std_logic_vector(14 downto 0);
  signal pgassign124 : std_logic_vector(31 downto 0);
  signal pgassign125 : std_logic_vector(31 downto 0);
  signal pgassign126 : std_logic_vector(3 downto 0);
  signal pgassign127 : std_logic_vector(14 downto 0);
  signal pgassign128 : std_logic_vector(31 downto 0);
  signal pgassign129 : std_logic_vector(31 downto 0);
  signal pgassign130 : std_logic_vector(3 downto 0);
  signal pgassign131 : std_logic_vector(14 downto 0);
  signal pgassign132 : std_logic_vector(31 downto 0);
  signal pgassign133 : std_logic_vector(31 downto 0);
  signal pgassign134 : std_logic_vector(3 downto 0);
  signal pgassign135 : std_logic_vector(14 downto 0);
  signal pgassign136 : std_logic_vector(31 downto 0);
  signal pgassign137 : std_logic_vector(31 downto 0);
  signal pgassign138 : std_logic_vector(3 downto 0);
  signal pgassign139 : std_logic_vector(14 downto 0);
  signal pgassign140 : std_logic_vector(31 downto 0);
  signal pgassign141 : std_logic_vector(31 downto 0);
  signal pgassign142 : std_logic_vector(3 downto 0);
  signal pgassign143 : std_logic_vector(14 downto 0);
  signal pgassign144 : std_logic_vector(31 downto 0);
  signal pgassign145 : std_logic_vector(31 downto 0);
  signal pgassign146 : std_logic_vector(3 downto 0);
  signal pgassign147 : std_logic_vector(14 downto 0);
  signal pgassign148 : std_logic_vector(31 downto 0);
  signal pgassign149 : std_logic_vector(31 downto 0);
  signal pgassign150 : std_logic_vector(3 downto 0);
  signal pgassign151 : std_logic_vector(14 downto 0);
  signal pgassign152 : std_logic_vector(31 downto 0);
  signal pgassign153 : std_logic_vector(31 downto 0);
  signal pgassign154 : std_logic_vector(3 downto 0);
  signal pgassign155 : std_logic_vector(14 downto 0);
  signal pgassign156 : std_logic_vector(31 downto 0);
  signal pgassign157 : std_logic_vector(31 downto 0);
  signal pgassign158 : std_logic_vector(3 downto 0);
  signal pgassign159 : std_logic_vector(14 downto 0);
  signal pgassign160 : std_logic_vector(31 downto 0);
  signal pgassign161 : std_logic_vector(31 downto 0);
  signal pgassign162 : std_logic_vector(3 downto 0);
  signal pgassign163 : std_logic_vector(14 downto 0);
  signal pgassign164 : std_logic_vector(31 downto 0);
  signal pgassign165 : std_logic_vector(31 downto 0);
  signal pgassign166 : std_logic_vector(3 downto 0);
  signal pgassign167 : std_logic_vector(14 downto 0);
  signal pgassign168 : std_logic_vector(31 downto 0);
  signal pgassign169 : std_logic_vector(31 downto 0);
  signal pgassign170 : std_logic_vector(3 downto 0);
  signal pgassign171 : std_logic_vector(14 downto 0);
  signal pgassign172 : std_logic_vector(31 downto 0);
  signal pgassign173 : std_logic_vector(31 downto 0);
  signal pgassign174 : std_logic_vector(3 downto 0);
  signal pgassign175 : std_logic_vector(14 downto 0);
  signal pgassign176 : std_logic_vector(31 downto 0);
  signal pgassign177 : std_logic_vector(31 downto 0);
  signal pgassign178 : std_logic_vector(3 downto 0);
  signal pgassign179 : std_logic_vector(14 downto 0);
  signal pgassign180 : std_logic_vector(31 downto 0);
  signal pgassign181 : std_logic_vector(31 downto 0);
  signal pgassign182 : std_logic_vector(3 downto 0);
  signal pgassign183 : std_logic_vector(14 downto 0);
  signal pgassign184 : std_logic_vector(31 downto 0);
  signal pgassign185 : std_logic_vector(31 downto 0);
  signal pgassign186 : std_logic_vector(3 downto 0);
  signal pgassign187 : std_logic_vector(14 downto 0);
  signal pgassign188 : std_logic_vector(31 downto 0);
  signal pgassign189 : std_logic_vector(31 downto 0);
  signal pgassign190 : std_logic_vector(3 downto 0);
  signal pgassign191 : std_logic_vector(14 downto 0);
  signal pgassign192 : std_logic_vector(31 downto 0);
  signal pgassign193 : std_logic_vector(31 downto 0);
  signal pgassign194 : std_logic_vector(3 downto 0);
  signal pgassign195 : std_logic_vector(14 downto 0);
  signal pgassign196 : std_logic_vector(31 downto 0);
  signal pgassign197 : std_logic_vector(31 downto 0);
  signal pgassign198 : std_logic_vector(3 downto 0);
  signal pgassign199 : std_logic_vector(14 downto 0);
  signal pgassign200 : std_logic_vector(31 downto 0);
  signal pgassign201 : std_logic_vector(31 downto 0);
  signal pgassign202 : std_logic_vector(3 downto 0);
  signal pgassign203 : std_logic_vector(14 downto 0);
  signal pgassign204 : std_logic_vector(31 downto 0);
  signal pgassign205 : std_logic_vector(31 downto 0);
  signal pgassign206 : std_logic_vector(3 downto 0);
  signal pgassign207 : std_logic_vector(14 downto 0);
  signal pgassign208 : std_logic_vector(31 downto 0);
  signal pgassign209 : std_logic_vector(31 downto 0);
  signal pgassign210 : std_logic_vector(3 downto 0);
  signal pgassign211 : std_logic_vector(14 downto 0);
  signal pgassign212 : std_logic_vector(31 downto 0);
  signal pgassign213 : std_logic_vector(31 downto 0);
  signal pgassign214 : std_logic_vector(3 downto 0);
  signal pgassign215 : std_logic_vector(14 downto 0);
  signal pgassign216 : std_logic_vector(31 downto 0);
  signal pgassign217 : std_logic_vector(31 downto 0);
  signal pgassign218 : std_logic_vector(3 downto 0);
  signal pgassign219 : std_logic_vector(14 downto 0);
  signal pgassign220 : std_logic_vector(31 downto 0);
  signal pgassign221 : std_logic_vector(31 downto 0);
  signal pgassign222 : std_logic_vector(3 downto 0);
  signal pgassign223 : std_logic_vector(14 downto 0);
  signal pgassign224 : std_logic_vector(31 downto 0);
  signal pgassign225 : std_logic_vector(31 downto 0);
  signal pgassign226 : std_logic_vector(3 downto 0);
  signal pgassign227 : std_logic_vector(14 downto 0);
  signal pgassign228 : std_logic_vector(31 downto 0);
  signal pgassign229 : std_logic_vector(31 downto 0);
  signal pgassign230 : std_logic_vector(3 downto 0);
  signal pgassign231 : std_logic_vector(14 downto 0);
  signal pgassign232 : std_logic_vector(31 downto 0);
  signal pgassign233 : std_logic_vector(31 downto 0);
  signal pgassign234 : std_logic_vector(3 downto 0);
  signal pgassign235 : std_logic_vector(14 downto 0);
  signal pgassign236 : std_logic_vector(31 downto 0);
  signal pgassign237 : std_logic_vector(31 downto 0);
  signal pgassign238 : std_logic_vector(3 downto 0);
  signal pgassign239 : std_logic_vector(14 downto 0);
  signal pgassign240 : std_logic_vector(31 downto 0);
  signal pgassign241 : std_logic_vector(31 downto 0);
  signal pgassign242 : std_logic_vector(3 downto 0);
  signal pgassign243 : std_logic_vector(14 downto 0);
  signal pgassign244 : std_logic_vector(31 downto 0);
  signal pgassign245 : std_logic_vector(31 downto 0);
  signal pgassign246 : std_logic_vector(3 downto 0);
  signal pgassign247 : std_logic_vector(14 downto 0);
  signal pgassign248 : std_logic_vector(31 downto 0);
  signal pgassign249 : std_logic_vector(31 downto 0);
  signal pgassign250 : std_logic_vector(3 downto 0);
  signal pgassign251 : std_logic_vector(14 downto 0);
  signal pgassign252 : std_logic_vector(31 downto 0);
  signal pgassign253 : std_logic_vector(31 downto 0);
  signal pgassign254 : std_logic_vector(3 downto 0);
  signal pgassign255 : std_logic_vector(14 downto 0);
  signal pgassign256 : std_logic_vector(31 downto 0);
  signal pgassign257 : std_logic_vector(31 downto 0);
  signal pgassign258 : std_logic_vector(3 downto 0);
  signal pgassign259 : std_logic_vector(14 downto 0);
  signal pgassign260 : std_logic_vector(31 downto 0);
  signal pgassign261 : std_logic_vector(31 downto 0);
  signal pgassign262 : std_logic_vector(3 downto 0);
  signal pgassign263 : std_logic_vector(14 downto 0);
  signal pgassign264 : std_logic_vector(31 downto 0);
  signal pgassign265 : std_logic_vector(31 downto 0);
  signal pgassign266 : std_logic_vector(3 downto 0);
  signal pgassign267 : std_logic_vector(14 downto 0);
  signal pgassign268 : std_logic_vector(31 downto 0);
  signal pgassign269 : std_logic_vector(31 downto 0);
  signal pgassign270 : std_logic_vector(3 downto 0);
  signal pgassign271 : std_logic_vector(14 downto 0);
  signal pgassign272 : std_logic_vector(31 downto 0);
  signal pgassign273 : std_logic_vector(31 downto 0);
  signal pgassign274 : std_logic_vector(3 downto 0);
  signal pgassign275 : std_logic_vector(14 downto 0);
  signal pgassign276 : std_logic_vector(31 downto 0);
  signal pgassign277 : std_logic_vector(31 downto 0);
  signal pgassign278 : std_logic_vector(3 downto 0);
  signal pgassign279 : std_logic_vector(14 downto 0);
  signal pgassign280 : std_logic_vector(31 downto 0);
  signal pgassign281 : std_logic_vector(31 downto 0);
  signal pgassign282 : std_logic_vector(3 downto 0);
  signal pgassign283 : std_logic_vector(14 downto 0);
  signal pgassign284 : std_logic_vector(31 downto 0);
  signal pgassign285 : std_logic_vector(31 downto 0);
  signal pgassign286 : std_logic_vector(3 downto 0);
  signal pgassign287 : std_logic_vector(14 downto 0);
  signal pgassign288 : std_logic_vector(31 downto 0);
  signal pgassign289 : std_logic_vector(31 downto 0);
  signal pgassign290 : std_logic_vector(3 downto 0);
  signal pgassign291 : std_logic_vector(14 downto 0);
  signal pgassign292 : std_logic_vector(31 downto 0);
  signal pgassign293 : std_logic_vector(31 downto 0);
  signal pgassign294 : std_logic_vector(3 downto 0);
  signal pgassign295 : std_logic_vector(14 downto 0);
  signal pgassign296 : std_logic_vector(31 downto 0);
  signal pgassign297 : std_logic_vector(31 downto 0);
  signal pgassign298 : std_logic_vector(3 downto 0);
  signal pgassign299 : std_logic_vector(14 downto 0);
  signal pgassign300 : std_logic_vector(31 downto 0);
  signal pgassign301 : std_logic_vector(31 downto 0);
  signal pgassign302 : std_logic_vector(3 downto 0);
  signal pgassign303 : std_logic_vector(14 downto 0);
  signal pgassign304 : std_logic_vector(31 downto 0);
  signal pgassign305 : std_logic_vector(31 downto 0);
  signal pgassign306 : std_logic_vector(3 downto 0);
  signal pgassign307 : std_logic_vector(14 downto 0);
  signal pgassign308 : std_logic_vector(31 downto 0);
  signal pgassign309 : std_logic_vector(31 downto 0);
  signal pgassign310 : std_logic_vector(3 downto 0);
  signal pgassign311 : std_logic_vector(14 downto 0);
  signal pgassign312 : std_logic_vector(31 downto 0);
  signal pgassign313 : std_logic_vector(31 downto 0);
  signal pgassign314 : std_logic_vector(3 downto 0);
  signal pgassign315 : std_logic_vector(14 downto 0);
  signal pgassign316 : std_logic_vector(31 downto 0);
  signal pgassign317 : std_logic_vector(31 downto 0);
  signal pgassign318 : std_logic_vector(3 downto 0);
  signal pgassign319 : std_logic_vector(14 downto 0);
  signal pgassign320 : std_logic_vector(31 downto 0);
  signal pgassign321 : std_logic_vector(31 downto 0);
  signal pgassign322 : std_logic_vector(3 downto 0);
  signal pgassign323 : std_logic_vector(14 downto 0);
  signal pgassign324 : std_logic_vector(31 downto 0);
  signal pgassign325 : std_logic_vector(31 downto 0);
  signal pgassign326 : std_logic_vector(3 downto 0);
  signal pgassign327 : std_logic_vector(14 downto 0);
  signal pgassign328 : std_logic_vector(31 downto 0);
  signal pgassign329 : std_logic_vector(31 downto 0);
  signal pgassign330 : std_logic_vector(3 downto 0);
  signal pgassign331 : std_logic_vector(14 downto 0);
  signal pgassign332 : std_logic_vector(31 downto 0);
  signal pgassign333 : std_logic_vector(31 downto 0);
  signal pgassign334 : std_logic_vector(3 downto 0);
  signal pgassign335 : std_logic_vector(14 downto 0);
  signal pgassign336 : std_logic_vector(31 downto 0);
  signal pgassign337 : std_logic_vector(31 downto 0);
  signal pgassign338 : std_logic_vector(3 downto 0);
  signal pgassign339 : std_logic_vector(14 downto 0);
  signal pgassign340 : std_logic_vector(31 downto 0);
  signal pgassign341 : std_logic_vector(31 downto 0);
  signal pgassign342 : std_logic_vector(3 downto 0);
  signal pgassign343 : std_logic_vector(14 downto 0);
  signal pgassign344 : std_logic_vector(31 downto 0);
  signal pgassign345 : std_logic_vector(31 downto 0);
  signal pgassign346 : std_logic_vector(3 downto 0);
  signal pgassign347 : std_logic_vector(14 downto 0);
  signal pgassign348 : std_logic_vector(31 downto 0);
  signal pgassign349 : std_logic_vector(31 downto 0);
  signal pgassign350 : std_logic_vector(3 downto 0);
  signal pgassign351 : std_logic_vector(14 downto 0);
  signal pgassign352 : std_logic_vector(31 downto 0);
  signal pgassign353 : std_logic_vector(31 downto 0);
  signal pgassign354 : std_logic_vector(3 downto 0);
  signal pgassign355 : std_logic_vector(14 downto 0);
  signal pgassign356 : std_logic_vector(31 downto 0);
  signal pgassign357 : std_logic_vector(31 downto 0);
  signal pgassign358 : std_logic_vector(3 downto 0);
  signal pgassign359 : std_logic_vector(14 downto 0);
  signal pgassign360 : std_logic_vector(31 downto 0);
  signal pgassign361 : std_logic_vector(31 downto 0);
  signal pgassign362 : std_logic_vector(3 downto 0);
  signal pgassign363 : std_logic_vector(14 downto 0);
  signal pgassign364 : std_logic_vector(31 downto 0);
  signal pgassign365 : std_logic_vector(31 downto 0);
  signal pgassign366 : std_logic_vector(3 downto 0);
  signal pgassign367 : std_logic_vector(14 downto 0);
  signal pgassign368 : std_logic_vector(31 downto 0);
  signal pgassign369 : std_logic_vector(31 downto 0);
  signal pgassign370 : std_logic_vector(3 downto 0);
  signal pgassign371 : std_logic_vector(14 downto 0);
  signal pgassign372 : std_logic_vector(31 downto 0);
  signal pgassign373 : std_logic_vector(31 downto 0);
  signal pgassign374 : std_logic_vector(3 downto 0);
  signal pgassign375 : std_logic_vector(14 downto 0);
  signal pgassign376 : std_logic_vector(31 downto 0);
  signal pgassign377 : std_logic_vector(31 downto 0);
  signal pgassign378 : std_logic_vector(3 downto 0);
  signal pgassign379 : std_logic_vector(14 downto 0);
  signal pgassign380 : std_logic_vector(31 downto 0);
  signal pgassign381 : std_logic_vector(31 downto 0);
  signal pgassign382 : std_logic_vector(3 downto 0);
  signal pgassign383 : std_logic_vector(14 downto 0);
  signal pgassign384 : std_logic_vector(31 downto 0);
  signal pgassign385 : std_logic_vector(31 downto 0);
  signal pgassign386 : std_logic_vector(3 downto 0);
  signal pgassign387 : std_logic_vector(14 downto 0);
  signal pgassign388 : std_logic_vector(31 downto 0);
  signal pgassign389 : std_logic_vector(31 downto 0);
  signal pgassign390 : std_logic_vector(3 downto 0);
  signal pgassign391 : std_logic_vector(14 downto 0);
  signal pgassign392 : std_logic_vector(31 downto 0);
  signal pgassign393 : std_logic_vector(31 downto 0);
  signal pgassign394 : std_logic_vector(3 downto 0);
  signal pgassign395 : std_logic_vector(14 downto 0);
  signal pgassign396 : std_logic_vector(31 downto 0);
  signal pgassign397 : std_logic_vector(31 downto 0);
  signal pgassign398 : std_logic_vector(3 downto 0);
  signal pgassign399 : std_logic_vector(14 downto 0);
  signal pgassign400 : std_logic_vector(31 downto 0);
  signal pgassign401 : std_logic_vector(31 downto 0);
  signal pgassign402 : std_logic_vector(3 downto 0);
  signal pgassign403 : std_logic_vector(14 downto 0);
  signal pgassign404 : std_logic_vector(31 downto 0);
  signal pgassign405 : std_logic_vector(31 downto 0);
  signal pgassign406 : std_logic_vector(3 downto 0);
  signal pgassign407 : std_logic_vector(14 downto 0);
  signal pgassign408 : std_logic_vector(31 downto 0);
  signal pgassign409 : std_logic_vector(31 downto 0);
  signal pgassign410 : std_logic_vector(3 downto 0);
  signal pgassign411 : std_logic_vector(14 downto 0);
  signal pgassign412 : std_logic_vector(31 downto 0);
  signal pgassign413 : std_logic_vector(31 downto 0);
  signal pgassign414 : std_logic_vector(3 downto 0);
  signal pgassign415 : std_logic_vector(14 downto 0);
  signal pgassign416 : std_logic_vector(31 downto 0);
  signal pgassign417 : std_logic_vector(31 downto 0);
  signal pgassign418 : std_logic_vector(3 downto 0);
  signal pgassign419 : std_logic_vector(14 downto 0);
  signal pgassign420 : std_logic_vector(31 downto 0);
  signal pgassign421 : std_logic_vector(31 downto 0);
  signal pgassign422 : std_logic_vector(3 downto 0);
  signal pgassign423 : std_logic_vector(14 downto 0);
  signal pgassign424 : std_logic_vector(31 downto 0);
  signal pgassign425 : std_logic_vector(31 downto 0);
  signal pgassign426 : std_logic_vector(3 downto 0);
  signal pgassign427 : std_logic_vector(14 downto 0);
  signal pgassign428 : std_logic_vector(31 downto 0);
  signal pgassign429 : std_logic_vector(31 downto 0);
  signal pgassign430 : std_logic_vector(3 downto 0);
  signal pgassign431 : std_logic_vector(14 downto 0);
  signal pgassign432 : std_logic_vector(31 downto 0);
  signal pgassign433 : std_logic_vector(31 downto 0);
  signal pgassign434 : std_logic_vector(3 downto 0);
  signal pgassign435 : std_logic_vector(14 downto 0);
  signal pgassign436 : std_logic_vector(31 downto 0);
  signal pgassign437 : std_logic_vector(31 downto 0);
  signal pgassign438 : std_logic_vector(3 downto 0);
  signal pgassign439 : std_logic_vector(14 downto 0);
  signal pgassign440 : std_logic_vector(31 downto 0);
  signal pgassign441 : std_logic_vector(31 downto 0);
  signal pgassign442 : std_logic_vector(3 downto 0);
  signal pgassign443 : std_logic_vector(14 downto 0);
  signal pgassign444 : std_logic_vector(31 downto 0);
  signal pgassign445 : std_logic_vector(31 downto 0);
  signal pgassign446 : std_logic_vector(3 downto 0);
  signal pgassign447 : std_logic_vector(14 downto 0);
  signal pgassign448 : std_logic_vector(31 downto 0);
  signal pgassign449 : std_logic_vector(31 downto 0);
  signal pgassign450 : std_logic_vector(3 downto 0);
  signal pgassign451 : std_logic_vector(14 downto 0);
  signal pgassign452 : std_logic_vector(31 downto 0);
  signal pgassign453 : std_logic_vector(31 downto 0);
  signal pgassign454 : std_logic_vector(3 downto 0);
  signal pgassign455 : std_logic_vector(14 downto 0);
  signal pgassign456 : std_logic_vector(31 downto 0);
  signal pgassign457 : std_logic_vector(31 downto 0);
  signal pgassign458 : std_logic_vector(3 downto 0);
  signal pgassign459 : std_logic_vector(14 downto 0);
  signal pgassign460 : std_logic_vector(31 downto 0);
  signal pgassign461 : std_logic_vector(31 downto 0);
  signal pgassign462 : std_logic_vector(3 downto 0);
  signal pgassign463 : std_logic_vector(14 downto 0);
  signal pgassign464 : std_logic_vector(31 downto 0);
  signal pgassign465 : std_logic_vector(31 downto 0);
  signal pgassign466 : std_logic_vector(3 downto 0);
  signal pgassign467 : std_logic_vector(14 downto 0);
  signal pgassign468 : std_logic_vector(31 downto 0);
  signal pgassign469 : std_logic_vector(31 downto 0);
  signal pgassign470 : std_logic_vector(3 downto 0);
  signal pgassign471 : std_logic_vector(14 downto 0);
  signal pgassign472 : std_logic_vector(31 downto 0);
  signal pgassign473 : std_logic_vector(31 downto 0);
  signal pgassign474 : std_logic_vector(3 downto 0);
  signal pgassign475 : std_logic_vector(14 downto 0);
  signal pgassign476 : std_logic_vector(31 downto 0);
  signal pgassign477 : std_logic_vector(31 downto 0);
  signal pgassign478 : std_logic_vector(3 downto 0);
  signal pgassign479 : std_logic_vector(14 downto 0);
  signal pgassign480 : std_logic_vector(31 downto 0);
  signal pgassign481 : std_logic_vector(31 downto 0);
  signal pgassign482 : std_logic_vector(3 downto 0);
  signal pgassign483 : std_logic_vector(14 downto 0);
  signal pgassign484 : std_logic_vector(31 downto 0);
  signal pgassign485 : std_logic_vector(31 downto 0);
  signal pgassign486 : std_logic_vector(3 downto 0);
  signal pgassign487 : std_logic_vector(14 downto 0);
  signal pgassign488 : std_logic_vector(31 downto 0);
  signal pgassign489 : std_logic_vector(31 downto 0);
  signal pgassign490 : std_logic_vector(3 downto 0);
  signal pgassign491 : std_logic_vector(14 downto 0);
  signal pgassign492 : std_logic_vector(31 downto 0);
  signal pgassign493 : std_logic_vector(31 downto 0);
  signal pgassign494 : std_logic_vector(3 downto 0);
  signal pgassign495 : std_logic_vector(14 downto 0);
  signal pgassign496 : std_logic_vector(31 downto 0);
  signal pgassign497 : std_logic_vector(31 downto 0);
  signal pgassign498 : std_logic_vector(3 downto 0);
  signal pgassign499 : std_logic_vector(14 downto 0);
  signal pgassign500 : std_logic_vector(31 downto 0);
  signal pgassign501 : std_logic_vector(31 downto 0);
  signal pgassign502 : std_logic_vector(3 downto 0);
  signal pgassign503 : std_logic_vector(14 downto 0);
  signal pgassign504 : std_logic_vector(31 downto 0);
  signal pgassign505 : std_logic_vector(31 downto 0);
  signal pgassign506 : std_logic_vector(3 downto 0);
  signal pgassign507 : std_logic_vector(14 downto 0);
  signal pgassign508 : std_logic_vector(31 downto 0);
  signal pgassign509 : std_logic_vector(31 downto 0);
  signal pgassign510 : std_logic_vector(3 downto 0);
  signal pgassign511 : std_logic_vector(14 downto 0);
  signal pgassign512 : std_logic_vector(31 downto 0);
  signal pgassign513 : std_logic_vector(31 downto 0);
  signal pgassign514 : std_logic_vector(3 downto 0);

begin

  -- Internal assignments

  pgassign1(0 to 0) <= B"1";
  pgassign2(0 to 30) <= B"0000000000000000000000000000000";
  pgassign3(14 downto 14) <= B"1";
  pgassign3(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign4(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign4(0 downto 0) <= BRAM_Dout_A(0 to 0);
  BRAM_Din_A(0 to 0) <= pgassign5(0 downto 0);
  pgassign6(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign6(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign6(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign6(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign7(14 downto 14) <= B"1";
  pgassign7(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign8(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign8(0 downto 0) <= BRAM_Dout_B(0 to 0);
  BRAM_Din_B(0 to 0) <= pgassign9(0 downto 0);
  pgassign10(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign10(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign10(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign10(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign11(14 downto 14) <= B"1";
  pgassign11(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign12(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign12(0 downto 0) <= BRAM_Dout_A(1 to 1);
  BRAM_Din_A(1 to 1) <= pgassign13(0 downto 0);
  pgassign14(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign14(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign14(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign14(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign15(14 downto 14) <= B"1";
  pgassign15(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign16(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign16(0 downto 0) <= BRAM_Dout_B(1 to 1);
  BRAM_Din_B(1 to 1) <= pgassign17(0 downto 0);
  pgassign18(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign18(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign18(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign18(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign19(14 downto 14) <= B"1";
  pgassign19(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign20(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign20(0 downto 0) <= BRAM_Dout_A(2 to 2);
  BRAM_Din_A(2 to 2) <= pgassign21(0 downto 0);
  pgassign22(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign22(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign22(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign22(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign23(14 downto 14) <= B"1";
  pgassign23(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign24(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign24(0 downto 0) <= BRAM_Dout_B(2 to 2);
  BRAM_Din_B(2 to 2) <= pgassign25(0 downto 0);
  pgassign26(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign26(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign26(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign26(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign27(14 downto 14) <= B"1";
  pgassign27(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign28(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign28(0 downto 0) <= BRAM_Dout_A(3 to 3);
  BRAM_Din_A(3 to 3) <= pgassign29(0 downto 0);
  pgassign30(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign30(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign30(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign30(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign31(14 downto 14) <= B"1";
  pgassign31(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign32(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign32(0 downto 0) <= BRAM_Dout_B(3 to 3);
  BRAM_Din_B(3 to 3) <= pgassign33(0 downto 0);
  pgassign34(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign34(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign34(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign34(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign35(14 downto 14) <= B"1";
  pgassign35(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign36(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign36(0 downto 0) <= BRAM_Dout_A(4 to 4);
  BRAM_Din_A(4 to 4) <= pgassign37(0 downto 0);
  pgassign38(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign38(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign38(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign38(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign39(14 downto 14) <= B"1";
  pgassign39(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign40(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign40(0 downto 0) <= BRAM_Dout_B(4 to 4);
  BRAM_Din_B(4 to 4) <= pgassign41(0 downto 0);
  pgassign42(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign42(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign42(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign42(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign43(14 downto 14) <= B"1";
  pgassign43(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign44(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign44(0 downto 0) <= BRAM_Dout_A(5 to 5);
  BRAM_Din_A(5 to 5) <= pgassign45(0 downto 0);
  pgassign46(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign46(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign46(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign46(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign47(14 downto 14) <= B"1";
  pgassign47(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign48(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign48(0 downto 0) <= BRAM_Dout_B(5 to 5);
  BRAM_Din_B(5 to 5) <= pgassign49(0 downto 0);
  pgassign50(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign50(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign50(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign50(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign51(14 downto 14) <= B"1";
  pgassign51(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign52(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign52(0 downto 0) <= BRAM_Dout_A(6 to 6);
  BRAM_Din_A(6 to 6) <= pgassign53(0 downto 0);
  pgassign54(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign54(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign54(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign54(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign55(14 downto 14) <= B"1";
  pgassign55(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign56(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign56(0 downto 0) <= BRAM_Dout_B(6 to 6);
  BRAM_Din_B(6 to 6) <= pgassign57(0 downto 0);
  pgassign58(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign58(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign58(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign58(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign59(14 downto 14) <= B"1";
  pgassign59(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign60(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign60(0 downto 0) <= BRAM_Dout_A(7 to 7);
  BRAM_Din_A(7 to 7) <= pgassign61(0 downto 0);
  pgassign62(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign62(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign62(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign62(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign63(14 downto 14) <= B"1";
  pgassign63(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign64(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign64(0 downto 0) <= BRAM_Dout_B(7 to 7);
  BRAM_Din_B(7 to 7) <= pgassign65(0 downto 0);
  pgassign66(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign66(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign66(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign66(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign67(14 downto 14) <= B"1";
  pgassign67(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign68(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign68(0 downto 0) <= BRAM_Dout_A(8 to 8);
  BRAM_Din_A(8 to 8) <= pgassign69(0 downto 0);
  pgassign70(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign70(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign70(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign70(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign71(14 downto 14) <= B"1";
  pgassign71(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign72(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign72(0 downto 0) <= BRAM_Dout_B(8 to 8);
  BRAM_Din_B(8 to 8) <= pgassign73(0 downto 0);
  pgassign74(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign74(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign74(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign74(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign75(14 downto 14) <= B"1";
  pgassign75(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign76(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign76(0 downto 0) <= BRAM_Dout_A(9 to 9);
  BRAM_Din_A(9 to 9) <= pgassign77(0 downto 0);
  pgassign78(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign78(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign78(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign78(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign79(14 downto 14) <= B"1";
  pgassign79(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign80(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign80(0 downto 0) <= BRAM_Dout_B(9 to 9);
  BRAM_Din_B(9 to 9) <= pgassign81(0 downto 0);
  pgassign82(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign82(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign82(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign82(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign83(14 downto 14) <= B"1";
  pgassign83(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign84(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign84(0 downto 0) <= BRAM_Dout_A(10 to 10);
  BRAM_Din_A(10 to 10) <= pgassign85(0 downto 0);
  pgassign86(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign86(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign86(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign86(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign87(14 downto 14) <= B"1";
  pgassign87(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign88(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign88(0 downto 0) <= BRAM_Dout_B(10 to 10);
  BRAM_Din_B(10 to 10) <= pgassign89(0 downto 0);
  pgassign90(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign90(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign90(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign90(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign91(14 downto 14) <= B"1";
  pgassign91(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign92(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign92(0 downto 0) <= BRAM_Dout_A(11 to 11);
  BRAM_Din_A(11 to 11) <= pgassign93(0 downto 0);
  pgassign94(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign94(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign94(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign94(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign95(14 downto 14) <= B"1";
  pgassign95(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign96(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign96(0 downto 0) <= BRAM_Dout_B(11 to 11);
  BRAM_Din_B(11 to 11) <= pgassign97(0 downto 0);
  pgassign98(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign98(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign98(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign98(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign99(14 downto 14) <= B"1";
  pgassign99(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign100(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign100(0 downto 0) <= BRAM_Dout_A(12 to 12);
  BRAM_Din_A(12 to 12) <= pgassign101(0 downto 0);
  pgassign102(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign102(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign102(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign102(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign103(14 downto 14) <= B"1";
  pgassign103(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign104(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign104(0 downto 0) <= BRAM_Dout_B(12 to 12);
  BRAM_Din_B(12 to 12) <= pgassign105(0 downto 0);
  pgassign106(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign106(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign106(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign106(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign107(14 downto 14) <= B"1";
  pgassign107(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign108(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign108(0 downto 0) <= BRAM_Dout_A(13 to 13);
  BRAM_Din_A(13 to 13) <= pgassign109(0 downto 0);
  pgassign110(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign110(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign110(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign110(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign111(14 downto 14) <= B"1";
  pgassign111(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign112(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign112(0 downto 0) <= BRAM_Dout_B(13 to 13);
  BRAM_Din_B(13 to 13) <= pgassign113(0 downto 0);
  pgassign114(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign114(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign114(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign114(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign115(14 downto 14) <= B"1";
  pgassign115(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign116(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign116(0 downto 0) <= BRAM_Dout_A(14 to 14);
  BRAM_Din_A(14 to 14) <= pgassign117(0 downto 0);
  pgassign118(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign118(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign118(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign118(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign119(14 downto 14) <= B"1";
  pgassign119(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign120(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign120(0 downto 0) <= BRAM_Dout_B(14 to 14);
  BRAM_Din_B(14 to 14) <= pgassign121(0 downto 0);
  pgassign122(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign122(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign122(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign122(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign123(14 downto 14) <= B"1";
  pgassign123(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign124(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign124(0 downto 0) <= BRAM_Dout_A(15 to 15);
  BRAM_Din_A(15 to 15) <= pgassign125(0 downto 0);
  pgassign126(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign126(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign126(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign126(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign127(14 downto 14) <= B"1";
  pgassign127(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign128(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign128(0 downto 0) <= BRAM_Dout_B(15 to 15);
  BRAM_Din_B(15 to 15) <= pgassign129(0 downto 0);
  pgassign130(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign130(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign130(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign130(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign131(14 downto 14) <= B"1";
  pgassign131(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign132(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign132(0 downto 0) <= BRAM_Dout_A(16 to 16);
  BRAM_Din_A(16 to 16) <= pgassign133(0 downto 0);
  pgassign134(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign134(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign134(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign134(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign135(14 downto 14) <= B"1";
  pgassign135(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign136(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign136(0 downto 0) <= BRAM_Dout_B(16 to 16);
  BRAM_Din_B(16 to 16) <= pgassign137(0 downto 0);
  pgassign138(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign138(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign138(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign138(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign139(14 downto 14) <= B"1";
  pgassign139(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign140(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign140(0 downto 0) <= BRAM_Dout_A(17 to 17);
  BRAM_Din_A(17 to 17) <= pgassign141(0 downto 0);
  pgassign142(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign142(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign142(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign142(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign143(14 downto 14) <= B"1";
  pgassign143(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign144(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign144(0 downto 0) <= BRAM_Dout_B(17 to 17);
  BRAM_Din_B(17 to 17) <= pgassign145(0 downto 0);
  pgassign146(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign146(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign146(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign146(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign147(14 downto 14) <= B"1";
  pgassign147(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign148(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign148(0 downto 0) <= BRAM_Dout_A(18 to 18);
  BRAM_Din_A(18 to 18) <= pgassign149(0 downto 0);
  pgassign150(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign150(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign150(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign150(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign151(14 downto 14) <= B"1";
  pgassign151(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign152(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign152(0 downto 0) <= BRAM_Dout_B(18 to 18);
  BRAM_Din_B(18 to 18) <= pgassign153(0 downto 0);
  pgassign154(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign154(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign154(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign154(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign155(14 downto 14) <= B"1";
  pgassign155(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign156(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign156(0 downto 0) <= BRAM_Dout_A(19 to 19);
  BRAM_Din_A(19 to 19) <= pgassign157(0 downto 0);
  pgassign158(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign158(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign158(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign158(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign159(14 downto 14) <= B"1";
  pgassign159(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign160(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign160(0 downto 0) <= BRAM_Dout_B(19 to 19);
  BRAM_Din_B(19 to 19) <= pgassign161(0 downto 0);
  pgassign162(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign162(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign162(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign162(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign163(14 downto 14) <= B"1";
  pgassign163(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign164(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign164(0 downto 0) <= BRAM_Dout_A(20 to 20);
  BRAM_Din_A(20 to 20) <= pgassign165(0 downto 0);
  pgassign166(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign166(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign166(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign166(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign167(14 downto 14) <= B"1";
  pgassign167(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign168(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign168(0 downto 0) <= BRAM_Dout_B(20 to 20);
  BRAM_Din_B(20 to 20) <= pgassign169(0 downto 0);
  pgassign170(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign170(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign170(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign170(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign171(14 downto 14) <= B"1";
  pgassign171(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign172(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign172(0 downto 0) <= BRAM_Dout_A(21 to 21);
  BRAM_Din_A(21 to 21) <= pgassign173(0 downto 0);
  pgassign174(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign174(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign174(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign174(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign175(14 downto 14) <= B"1";
  pgassign175(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign176(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign176(0 downto 0) <= BRAM_Dout_B(21 to 21);
  BRAM_Din_B(21 to 21) <= pgassign177(0 downto 0);
  pgassign178(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign178(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign178(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign178(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign179(14 downto 14) <= B"1";
  pgassign179(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign180(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign180(0 downto 0) <= BRAM_Dout_A(22 to 22);
  BRAM_Din_A(22 to 22) <= pgassign181(0 downto 0);
  pgassign182(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign182(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign182(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign182(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign183(14 downto 14) <= B"1";
  pgassign183(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign184(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign184(0 downto 0) <= BRAM_Dout_B(22 to 22);
  BRAM_Din_B(22 to 22) <= pgassign185(0 downto 0);
  pgassign186(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign186(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign186(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign186(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign187(14 downto 14) <= B"1";
  pgassign187(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign188(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign188(0 downto 0) <= BRAM_Dout_A(23 to 23);
  BRAM_Din_A(23 to 23) <= pgassign189(0 downto 0);
  pgassign190(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign190(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign190(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign190(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign191(14 downto 14) <= B"1";
  pgassign191(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign192(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign192(0 downto 0) <= BRAM_Dout_B(23 to 23);
  BRAM_Din_B(23 to 23) <= pgassign193(0 downto 0);
  pgassign194(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign194(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign194(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign194(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign195(14 downto 14) <= B"1";
  pgassign195(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign196(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign196(0 downto 0) <= BRAM_Dout_A(24 to 24);
  BRAM_Din_A(24 to 24) <= pgassign197(0 downto 0);
  pgassign198(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign198(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign198(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign198(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign199(14 downto 14) <= B"1";
  pgassign199(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign200(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign200(0 downto 0) <= BRAM_Dout_B(24 to 24);
  BRAM_Din_B(24 to 24) <= pgassign201(0 downto 0);
  pgassign202(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign202(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign202(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign202(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign203(14 downto 14) <= B"1";
  pgassign203(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign204(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign204(0 downto 0) <= BRAM_Dout_A(25 to 25);
  BRAM_Din_A(25 to 25) <= pgassign205(0 downto 0);
  pgassign206(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign206(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign206(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign206(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign207(14 downto 14) <= B"1";
  pgassign207(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign208(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign208(0 downto 0) <= BRAM_Dout_B(25 to 25);
  BRAM_Din_B(25 to 25) <= pgassign209(0 downto 0);
  pgassign210(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign210(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign210(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign210(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign211(14 downto 14) <= B"1";
  pgassign211(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign212(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign212(0 downto 0) <= BRAM_Dout_A(26 to 26);
  BRAM_Din_A(26 to 26) <= pgassign213(0 downto 0);
  pgassign214(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign214(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign214(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign214(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign215(14 downto 14) <= B"1";
  pgassign215(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign216(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign216(0 downto 0) <= BRAM_Dout_B(26 to 26);
  BRAM_Din_B(26 to 26) <= pgassign217(0 downto 0);
  pgassign218(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign218(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign218(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign218(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign219(14 downto 14) <= B"1";
  pgassign219(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign220(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign220(0 downto 0) <= BRAM_Dout_A(27 to 27);
  BRAM_Din_A(27 to 27) <= pgassign221(0 downto 0);
  pgassign222(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign222(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign222(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign222(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign223(14 downto 14) <= B"1";
  pgassign223(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign224(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign224(0 downto 0) <= BRAM_Dout_B(27 to 27);
  BRAM_Din_B(27 to 27) <= pgassign225(0 downto 0);
  pgassign226(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign226(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign226(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign226(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign227(14 downto 14) <= B"1";
  pgassign227(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign228(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign228(0 downto 0) <= BRAM_Dout_A(28 to 28);
  BRAM_Din_A(28 to 28) <= pgassign229(0 downto 0);
  pgassign230(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign230(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign230(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign230(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign231(14 downto 14) <= B"1";
  pgassign231(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign232(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign232(0 downto 0) <= BRAM_Dout_B(28 to 28);
  BRAM_Din_B(28 to 28) <= pgassign233(0 downto 0);
  pgassign234(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign234(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign234(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign234(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign235(14 downto 14) <= B"1";
  pgassign235(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign236(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign236(0 downto 0) <= BRAM_Dout_A(29 to 29);
  BRAM_Din_A(29 to 29) <= pgassign237(0 downto 0);
  pgassign238(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign238(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign238(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign238(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign239(14 downto 14) <= B"1";
  pgassign239(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign240(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign240(0 downto 0) <= BRAM_Dout_B(29 to 29);
  BRAM_Din_B(29 to 29) <= pgassign241(0 downto 0);
  pgassign242(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign242(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign242(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign242(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign243(14 downto 14) <= B"1";
  pgassign243(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign244(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign244(0 downto 0) <= BRAM_Dout_A(30 to 30);
  BRAM_Din_A(30 to 30) <= pgassign245(0 downto 0);
  pgassign246(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign246(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign246(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign246(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign247(14 downto 14) <= B"1";
  pgassign247(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign248(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign248(0 downto 0) <= BRAM_Dout_B(30 to 30);
  BRAM_Din_B(30 to 30) <= pgassign249(0 downto 0);
  pgassign250(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign250(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign250(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign250(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign251(14 downto 14) <= B"1";
  pgassign251(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign252(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign252(0 downto 0) <= BRAM_Dout_A(31 to 31);
  BRAM_Din_A(31 to 31) <= pgassign253(0 downto 0);
  pgassign254(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign254(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign254(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign254(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign255(14 downto 14) <= B"1";
  pgassign255(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign256(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign256(0 downto 0) <= BRAM_Dout_B(31 to 31);
  BRAM_Din_B(31 to 31) <= pgassign257(0 downto 0);
  pgassign258(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign258(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign258(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign258(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign259(14 downto 14) <= B"1";
  pgassign259(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign260(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign260(0 downto 0) <= BRAM_Dout_A(32 to 32);
  BRAM_Din_A(32 to 32) <= pgassign261(0 downto 0);
  pgassign262(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign262(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign262(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign262(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign263(14 downto 14) <= B"1";
  pgassign263(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign264(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign264(0 downto 0) <= BRAM_Dout_B(32 to 32);
  BRAM_Din_B(32 to 32) <= pgassign265(0 downto 0);
  pgassign266(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign266(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign266(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign266(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign267(14 downto 14) <= B"1";
  pgassign267(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign268(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign268(0 downto 0) <= BRAM_Dout_A(33 to 33);
  BRAM_Din_A(33 to 33) <= pgassign269(0 downto 0);
  pgassign270(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign270(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign270(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign270(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign271(14 downto 14) <= B"1";
  pgassign271(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign272(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign272(0 downto 0) <= BRAM_Dout_B(33 to 33);
  BRAM_Din_B(33 to 33) <= pgassign273(0 downto 0);
  pgassign274(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign274(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign274(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign274(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign275(14 downto 14) <= B"1";
  pgassign275(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign276(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign276(0 downto 0) <= BRAM_Dout_A(34 to 34);
  BRAM_Din_A(34 to 34) <= pgassign277(0 downto 0);
  pgassign278(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign278(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign278(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign278(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign279(14 downto 14) <= B"1";
  pgassign279(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign280(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign280(0 downto 0) <= BRAM_Dout_B(34 to 34);
  BRAM_Din_B(34 to 34) <= pgassign281(0 downto 0);
  pgassign282(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign282(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign282(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign282(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign283(14 downto 14) <= B"1";
  pgassign283(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign284(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign284(0 downto 0) <= BRAM_Dout_A(35 to 35);
  BRAM_Din_A(35 to 35) <= pgassign285(0 downto 0);
  pgassign286(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign286(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign286(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign286(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign287(14 downto 14) <= B"1";
  pgassign287(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign288(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign288(0 downto 0) <= BRAM_Dout_B(35 to 35);
  BRAM_Din_B(35 to 35) <= pgassign289(0 downto 0);
  pgassign290(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign290(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign290(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign290(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign291(14 downto 14) <= B"1";
  pgassign291(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign292(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign292(0 downto 0) <= BRAM_Dout_A(36 to 36);
  BRAM_Din_A(36 to 36) <= pgassign293(0 downto 0);
  pgassign294(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign294(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign294(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign294(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign295(14 downto 14) <= B"1";
  pgassign295(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign296(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign296(0 downto 0) <= BRAM_Dout_B(36 to 36);
  BRAM_Din_B(36 to 36) <= pgassign297(0 downto 0);
  pgassign298(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign298(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign298(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign298(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign299(14 downto 14) <= B"1";
  pgassign299(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign300(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign300(0 downto 0) <= BRAM_Dout_A(37 to 37);
  BRAM_Din_A(37 to 37) <= pgassign301(0 downto 0);
  pgassign302(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign302(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign302(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign302(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign303(14 downto 14) <= B"1";
  pgassign303(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign304(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign304(0 downto 0) <= BRAM_Dout_B(37 to 37);
  BRAM_Din_B(37 to 37) <= pgassign305(0 downto 0);
  pgassign306(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign306(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign306(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign306(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign307(14 downto 14) <= B"1";
  pgassign307(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign308(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign308(0 downto 0) <= BRAM_Dout_A(38 to 38);
  BRAM_Din_A(38 to 38) <= pgassign309(0 downto 0);
  pgassign310(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign310(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign310(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign310(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign311(14 downto 14) <= B"1";
  pgassign311(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign312(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign312(0 downto 0) <= BRAM_Dout_B(38 to 38);
  BRAM_Din_B(38 to 38) <= pgassign313(0 downto 0);
  pgassign314(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign314(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign314(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign314(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign315(14 downto 14) <= B"1";
  pgassign315(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign316(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign316(0 downto 0) <= BRAM_Dout_A(39 to 39);
  BRAM_Din_A(39 to 39) <= pgassign317(0 downto 0);
  pgassign318(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign318(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign318(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign318(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign319(14 downto 14) <= B"1";
  pgassign319(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign320(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign320(0 downto 0) <= BRAM_Dout_B(39 to 39);
  BRAM_Din_B(39 to 39) <= pgassign321(0 downto 0);
  pgassign322(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign322(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign322(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign322(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign323(14 downto 14) <= B"1";
  pgassign323(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign324(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign324(0 downto 0) <= BRAM_Dout_A(40 to 40);
  BRAM_Din_A(40 to 40) <= pgassign325(0 downto 0);
  pgassign326(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign326(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign326(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign326(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign327(14 downto 14) <= B"1";
  pgassign327(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign328(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign328(0 downto 0) <= BRAM_Dout_B(40 to 40);
  BRAM_Din_B(40 to 40) <= pgassign329(0 downto 0);
  pgassign330(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign330(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign330(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign330(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign331(14 downto 14) <= B"1";
  pgassign331(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign332(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign332(0 downto 0) <= BRAM_Dout_A(41 to 41);
  BRAM_Din_A(41 to 41) <= pgassign333(0 downto 0);
  pgassign334(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign334(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign334(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign334(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign335(14 downto 14) <= B"1";
  pgassign335(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign336(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign336(0 downto 0) <= BRAM_Dout_B(41 to 41);
  BRAM_Din_B(41 to 41) <= pgassign337(0 downto 0);
  pgassign338(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign338(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign338(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign338(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign339(14 downto 14) <= B"1";
  pgassign339(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign340(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign340(0 downto 0) <= BRAM_Dout_A(42 to 42);
  BRAM_Din_A(42 to 42) <= pgassign341(0 downto 0);
  pgassign342(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign342(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign342(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign342(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign343(14 downto 14) <= B"1";
  pgassign343(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign344(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign344(0 downto 0) <= BRAM_Dout_B(42 to 42);
  BRAM_Din_B(42 to 42) <= pgassign345(0 downto 0);
  pgassign346(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign346(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign346(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign346(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign347(14 downto 14) <= B"1";
  pgassign347(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign348(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign348(0 downto 0) <= BRAM_Dout_A(43 to 43);
  BRAM_Din_A(43 to 43) <= pgassign349(0 downto 0);
  pgassign350(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign350(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign350(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign350(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign351(14 downto 14) <= B"1";
  pgassign351(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign352(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign352(0 downto 0) <= BRAM_Dout_B(43 to 43);
  BRAM_Din_B(43 to 43) <= pgassign353(0 downto 0);
  pgassign354(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign354(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign354(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign354(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign355(14 downto 14) <= B"1";
  pgassign355(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign356(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign356(0 downto 0) <= BRAM_Dout_A(44 to 44);
  BRAM_Din_A(44 to 44) <= pgassign357(0 downto 0);
  pgassign358(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign358(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign358(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign358(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign359(14 downto 14) <= B"1";
  pgassign359(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign360(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign360(0 downto 0) <= BRAM_Dout_B(44 to 44);
  BRAM_Din_B(44 to 44) <= pgassign361(0 downto 0);
  pgassign362(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign362(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign362(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign362(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign363(14 downto 14) <= B"1";
  pgassign363(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign364(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign364(0 downto 0) <= BRAM_Dout_A(45 to 45);
  BRAM_Din_A(45 to 45) <= pgassign365(0 downto 0);
  pgassign366(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign366(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign366(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign366(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign367(14 downto 14) <= B"1";
  pgassign367(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign368(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign368(0 downto 0) <= BRAM_Dout_B(45 to 45);
  BRAM_Din_B(45 to 45) <= pgassign369(0 downto 0);
  pgassign370(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign370(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign370(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign370(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign371(14 downto 14) <= B"1";
  pgassign371(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign372(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign372(0 downto 0) <= BRAM_Dout_A(46 to 46);
  BRAM_Din_A(46 to 46) <= pgassign373(0 downto 0);
  pgassign374(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign374(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign374(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign374(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign375(14 downto 14) <= B"1";
  pgassign375(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign376(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign376(0 downto 0) <= BRAM_Dout_B(46 to 46);
  BRAM_Din_B(46 to 46) <= pgassign377(0 downto 0);
  pgassign378(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign378(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign378(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign378(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign379(14 downto 14) <= B"1";
  pgassign379(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign380(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign380(0 downto 0) <= BRAM_Dout_A(47 to 47);
  BRAM_Din_A(47 to 47) <= pgassign381(0 downto 0);
  pgassign382(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign382(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign382(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign382(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign383(14 downto 14) <= B"1";
  pgassign383(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign384(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign384(0 downto 0) <= BRAM_Dout_B(47 to 47);
  BRAM_Din_B(47 to 47) <= pgassign385(0 downto 0);
  pgassign386(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign386(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign386(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign386(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign387(14 downto 14) <= B"1";
  pgassign387(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign388(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign388(0 downto 0) <= BRAM_Dout_A(48 to 48);
  BRAM_Din_A(48 to 48) <= pgassign389(0 downto 0);
  pgassign390(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign390(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign390(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign390(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign391(14 downto 14) <= B"1";
  pgassign391(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign392(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign392(0 downto 0) <= BRAM_Dout_B(48 to 48);
  BRAM_Din_B(48 to 48) <= pgassign393(0 downto 0);
  pgassign394(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign394(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign394(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign394(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign395(14 downto 14) <= B"1";
  pgassign395(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign396(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign396(0 downto 0) <= BRAM_Dout_A(49 to 49);
  BRAM_Din_A(49 to 49) <= pgassign397(0 downto 0);
  pgassign398(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign398(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign398(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign398(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign399(14 downto 14) <= B"1";
  pgassign399(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign400(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign400(0 downto 0) <= BRAM_Dout_B(49 to 49);
  BRAM_Din_B(49 to 49) <= pgassign401(0 downto 0);
  pgassign402(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign402(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign402(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign402(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign403(14 downto 14) <= B"1";
  pgassign403(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign404(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign404(0 downto 0) <= BRAM_Dout_A(50 to 50);
  BRAM_Din_A(50 to 50) <= pgassign405(0 downto 0);
  pgassign406(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign406(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign406(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign406(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign407(14 downto 14) <= B"1";
  pgassign407(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign408(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign408(0 downto 0) <= BRAM_Dout_B(50 to 50);
  BRAM_Din_B(50 to 50) <= pgassign409(0 downto 0);
  pgassign410(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign410(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign410(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign410(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign411(14 downto 14) <= B"1";
  pgassign411(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign412(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign412(0 downto 0) <= BRAM_Dout_A(51 to 51);
  BRAM_Din_A(51 to 51) <= pgassign413(0 downto 0);
  pgassign414(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign414(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign414(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign414(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign415(14 downto 14) <= B"1";
  pgassign415(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign416(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign416(0 downto 0) <= BRAM_Dout_B(51 to 51);
  BRAM_Din_B(51 to 51) <= pgassign417(0 downto 0);
  pgassign418(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign418(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign418(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign418(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign419(14 downto 14) <= B"1";
  pgassign419(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign420(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign420(0 downto 0) <= BRAM_Dout_A(52 to 52);
  BRAM_Din_A(52 to 52) <= pgassign421(0 downto 0);
  pgassign422(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign422(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign422(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign422(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign423(14 downto 14) <= B"1";
  pgassign423(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign424(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign424(0 downto 0) <= BRAM_Dout_B(52 to 52);
  BRAM_Din_B(52 to 52) <= pgassign425(0 downto 0);
  pgassign426(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign426(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign426(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign426(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign427(14 downto 14) <= B"1";
  pgassign427(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign428(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign428(0 downto 0) <= BRAM_Dout_A(53 to 53);
  BRAM_Din_A(53 to 53) <= pgassign429(0 downto 0);
  pgassign430(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign430(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign430(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign430(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign431(14 downto 14) <= B"1";
  pgassign431(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign432(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign432(0 downto 0) <= BRAM_Dout_B(53 to 53);
  BRAM_Din_B(53 to 53) <= pgassign433(0 downto 0);
  pgassign434(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign434(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign434(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign434(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign435(14 downto 14) <= B"1";
  pgassign435(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign436(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign436(0 downto 0) <= BRAM_Dout_A(54 to 54);
  BRAM_Din_A(54 to 54) <= pgassign437(0 downto 0);
  pgassign438(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign438(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign438(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign438(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign439(14 downto 14) <= B"1";
  pgassign439(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign440(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign440(0 downto 0) <= BRAM_Dout_B(54 to 54);
  BRAM_Din_B(54 to 54) <= pgassign441(0 downto 0);
  pgassign442(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign442(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign442(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign442(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign443(14 downto 14) <= B"1";
  pgassign443(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign444(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign444(0 downto 0) <= BRAM_Dout_A(55 to 55);
  BRAM_Din_A(55 to 55) <= pgassign445(0 downto 0);
  pgassign446(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign446(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign446(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign446(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign447(14 downto 14) <= B"1";
  pgassign447(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign448(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign448(0 downto 0) <= BRAM_Dout_B(55 to 55);
  BRAM_Din_B(55 to 55) <= pgassign449(0 downto 0);
  pgassign450(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign450(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign450(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign450(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign451(14 downto 14) <= B"1";
  pgassign451(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign452(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign452(0 downto 0) <= BRAM_Dout_A(56 to 56);
  BRAM_Din_A(56 to 56) <= pgassign453(0 downto 0);
  pgassign454(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign454(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign454(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign454(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign455(14 downto 14) <= B"1";
  pgassign455(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign456(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign456(0 downto 0) <= BRAM_Dout_B(56 to 56);
  BRAM_Din_B(56 to 56) <= pgassign457(0 downto 0);
  pgassign458(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign458(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign458(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign458(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign459(14 downto 14) <= B"1";
  pgassign459(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign460(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign460(0 downto 0) <= BRAM_Dout_A(57 to 57);
  BRAM_Din_A(57 to 57) <= pgassign461(0 downto 0);
  pgassign462(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign462(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign462(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign462(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign463(14 downto 14) <= B"1";
  pgassign463(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign464(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign464(0 downto 0) <= BRAM_Dout_B(57 to 57);
  BRAM_Din_B(57 to 57) <= pgassign465(0 downto 0);
  pgassign466(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign466(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign466(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign466(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign467(14 downto 14) <= B"1";
  pgassign467(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign468(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign468(0 downto 0) <= BRAM_Dout_A(58 to 58);
  BRAM_Din_A(58 to 58) <= pgassign469(0 downto 0);
  pgassign470(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign470(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign470(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign470(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign471(14 downto 14) <= B"1";
  pgassign471(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign472(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign472(0 downto 0) <= BRAM_Dout_B(58 to 58);
  BRAM_Din_B(58 to 58) <= pgassign473(0 downto 0);
  pgassign474(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign474(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign474(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign474(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign475(14 downto 14) <= B"1";
  pgassign475(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign476(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign476(0 downto 0) <= BRAM_Dout_A(59 to 59);
  BRAM_Din_A(59 to 59) <= pgassign477(0 downto 0);
  pgassign478(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign478(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign478(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign478(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign479(14 downto 14) <= B"1";
  pgassign479(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign480(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign480(0 downto 0) <= BRAM_Dout_B(59 to 59);
  BRAM_Din_B(59 to 59) <= pgassign481(0 downto 0);
  pgassign482(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign482(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign482(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign482(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign483(14 downto 14) <= B"1";
  pgassign483(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign484(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign484(0 downto 0) <= BRAM_Dout_A(60 to 60);
  BRAM_Din_A(60 to 60) <= pgassign485(0 downto 0);
  pgassign486(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign486(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign486(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign486(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign487(14 downto 14) <= B"1";
  pgassign487(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign488(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign488(0 downto 0) <= BRAM_Dout_B(60 to 60);
  BRAM_Din_B(60 to 60) <= pgassign489(0 downto 0);
  pgassign490(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign490(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign490(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign490(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign491(14 downto 14) <= B"1";
  pgassign491(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign492(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign492(0 downto 0) <= BRAM_Dout_A(61 to 61);
  BRAM_Din_A(61 to 61) <= pgassign493(0 downto 0);
  pgassign494(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign494(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign494(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign494(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign495(14 downto 14) <= B"1";
  pgassign495(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign496(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign496(0 downto 0) <= BRAM_Dout_B(61 to 61);
  BRAM_Din_B(61 to 61) <= pgassign497(0 downto 0);
  pgassign498(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign498(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign498(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign498(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign499(14 downto 14) <= B"1";
  pgassign499(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign500(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign500(0 downto 0) <= BRAM_Dout_A(62 to 62);
  BRAM_Din_A(62 to 62) <= pgassign501(0 downto 0);
  pgassign502(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign502(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign502(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign502(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign503(14 downto 14) <= B"1";
  pgassign503(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign504(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign504(0 downto 0) <= BRAM_Dout_B(62 to 62);
  BRAM_Din_B(62 to 62) <= pgassign505(0 downto 0);
  pgassign506(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign506(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign506(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign506(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign507(14 downto 14) <= B"1";
  pgassign507(13 downto 0) <= BRAM_Addr_A(15 to 28);
  pgassign508(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign508(0 downto 0) <= BRAM_Dout_A(63 to 63);
  BRAM_Din_A(63 to 63) <= pgassign509(0 downto 0);
  pgassign510(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign510(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign510(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign510(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign511(14 downto 14) <= B"1";
  pgassign511(13 downto 0) <= BRAM_Addr_B(15 to 28);
  pgassign512(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign512(0 downto 0) <= BRAM_Dout_B(63 to 63);
  BRAM_Din_B(63 to 63) <= pgassign513(0 downto 0);
  pgassign514(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign514(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign514(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign514(0 downto 0) <= BRAM_WEN_B(7 to 7);
  net_gnd0 <= '0';
  net_gnd4(3 downto 0) <= B"0000";

  ramb16_0 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_0.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign3,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign4,
      DIPA => net_gnd4,
      DOA => pgassign5,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign6,
      ADDRB => pgassign7,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign8,
      DIPB => net_gnd4,
      DOB => pgassign9,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign10
    );

  ramb16_1 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_1.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign11,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign12,
      DIPA => net_gnd4,
      DOA => pgassign13,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign14,
      ADDRB => pgassign15,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign16,
      DIPB => net_gnd4,
      DOB => pgassign17,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign18
    );

  ramb16_2 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_2.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign19,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign20,
      DIPA => net_gnd4,
      DOA => pgassign21,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign22,
      ADDRB => pgassign23,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign24,
      DIPB => net_gnd4,
      DOB => pgassign25,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign26
    );

  ramb16_3 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_3.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign27,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign28,
      DIPA => net_gnd4,
      DOA => pgassign29,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign30,
      ADDRB => pgassign31,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign32,
      DIPB => net_gnd4,
      DOB => pgassign33,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign34
    );

  ramb16_4 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_4.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign35,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign36,
      DIPA => net_gnd4,
      DOA => pgassign37,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign38,
      ADDRB => pgassign39,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign40,
      DIPB => net_gnd4,
      DOB => pgassign41,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign42
    );

  ramb16_5 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_5.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign43,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign44,
      DIPA => net_gnd4,
      DOA => pgassign45,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign46,
      ADDRB => pgassign47,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign48,
      DIPB => net_gnd4,
      DOB => pgassign49,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign50
    );

  ramb16_6 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_6.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign51,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign52,
      DIPA => net_gnd4,
      DOA => pgassign53,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign54,
      ADDRB => pgassign55,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign56,
      DIPB => net_gnd4,
      DOB => pgassign57,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign58
    );

  ramb16_7 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_7.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign59,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign60,
      DIPA => net_gnd4,
      DOA => pgassign61,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign62,
      ADDRB => pgassign63,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign64,
      DIPB => net_gnd4,
      DOB => pgassign65,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign66
    );

  ramb16_8 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_8.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign67,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign68,
      DIPA => net_gnd4,
      DOA => pgassign69,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign70,
      ADDRB => pgassign71,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign72,
      DIPB => net_gnd4,
      DOB => pgassign73,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign74
    );

  ramb16_9 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_9.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign75,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign76,
      DIPA => net_gnd4,
      DOA => pgassign77,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign78,
      ADDRB => pgassign79,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign80,
      DIPB => net_gnd4,
      DOB => pgassign81,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign82
    );

  ramb16_10 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_10.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign83,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign84,
      DIPA => net_gnd4,
      DOA => pgassign85,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign86,
      ADDRB => pgassign87,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign88,
      DIPB => net_gnd4,
      DOB => pgassign89,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign90
    );

  ramb16_11 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_11.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign91,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign92,
      DIPA => net_gnd4,
      DOA => pgassign93,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign94,
      ADDRB => pgassign95,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign96,
      DIPB => net_gnd4,
      DOB => pgassign97,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign98
    );

  ramb16_12 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_12.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign99,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign100,
      DIPA => net_gnd4,
      DOA => pgassign101,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign102,
      ADDRB => pgassign103,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign104,
      DIPB => net_gnd4,
      DOB => pgassign105,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign106
    );

  ramb16_13 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_13.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign107,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign108,
      DIPA => net_gnd4,
      DOA => pgassign109,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign110,
      ADDRB => pgassign111,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign112,
      DIPB => net_gnd4,
      DOB => pgassign113,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign114
    );

  ramb16_14 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_14.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign115,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign116,
      DIPA => net_gnd4,
      DOA => pgassign117,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign118,
      ADDRB => pgassign119,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign120,
      DIPB => net_gnd4,
      DOB => pgassign121,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign122
    );

  ramb16_15 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_15.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign123,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign124,
      DIPA => net_gnd4,
      DOA => pgassign125,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign126,
      ADDRB => pgassign127,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign128,
      DIPB => net_gnd4,
      DOB => pgassign129,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign130
    );

  ramb16_16 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_16.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign131,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign132,
      DIPA => net_gnd4,
      DOA => pgassign133,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign134,
      ADDRB => pgassign135,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign136,
      DIPB => net_gnd4,
      DOB => pgassign137,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign138
    );

  ramb16_17 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_17.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign139,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign140,
      DIPA => net_gnd4,
      DOA => pgassign141,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign142,
      ADDRB => pgassign143,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign144,
      DIPB => net_gnd4,
      DOB => pgassign145,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign146
    );

  ramb16_18 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_18.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign147,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign148,
      DIPA => net_gnd4,
      DOA => pgassign149,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign150,
      ADDRB => pgassign151,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign152,
      DIPB => net_gnd4,
      DOB => pgassign153,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign154
    );

  ramb16_19 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_19.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign155,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign156,
      DIPA => net_gnd4,
      DOA => pgassign157,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign158,
      ADDRB => pgassign159,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign160,
      DIPB => net_gnd4,
      DOB => pgassign161,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign162
    );

  ramb16_20 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_20.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign163,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign164,
      DIPA => net_gnd4,
      DOA => pgassign165,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign166,
      ADDRB => pgassign167,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign168,
      DIPB => net_gnd4,
      DOB => pgassign169,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign170
    );

  ramb16_21 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_21.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign171,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign172,
      DIPA => net_gnd4,
      DOA => pgassign173,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign174,
      ADDRB => pgassign175,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign176,
      DIPB => net_gnd4,
      DOB => pgassign177,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign178
    );

  ramb16_22 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_22.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign179,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign180,
      DIPA => net_gnd4,
      DOA => pgassign181,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign182,
      ADDRB => pgassign183,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign184,
      DIPB => net_gnd4,
      DOB => pgassign185,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign186
    );

  ramb16_23 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_23.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign187,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign188,
      DIPA => net_gnd4,
      DOA => pgassign189,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign190,
      ADDRB => pgassign191,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign192,
      DIPB => net_gnd4,
      DOB => pgassign193,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign194
    );

  ramb16_24 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_24.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign195,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign196,
      DIPA => net_gnd4,
      DOA => pgassign197,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign198,
      ADDRB => pgassign199,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign200,
      DIPB => net_gnd4,
      DOB => pgassign201,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign202
    );

  ramb16_25 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_25.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign203,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign204,
      DIPA => net_gnd4,
      DOA => pgassign205,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign206,
      ADDRB => pgassign207,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign208,
      DIPB => net_gnd4,
      DOB => pgassign209,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign210
    );

  ramb16_26 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_26.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign211,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign212,
      DIPA => net_gnd4,
      DOA => pgassign213,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign214,
      ADDRB => pgassign215,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign216,
      DIPB => net_gnd4,
      DOB => pgassign217,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign218
    );

  ramb16_27 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_27.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign219,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign220,
      DIPA => net_gnd4,
      DOA => pgassign221,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign222,
      ADDRB => pgassign223,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign224,
      DIPB => net_gnd4,
      DOB => pgassign225,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign226
    );

  ramb16_28 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_28.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign227,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign228,
      DIPA => net_gnd4,
      DOA => pgassign229,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign230,
      ADDRB => pgassign231,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign232,
      DIPB => net_gnd4,
      DOB => pgassign233,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign234
    );

  ramb16_29 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_29.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign235,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign236,
      DIPA => net_gnd4,
      DOA => pgassign237,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign238,
      ADDRB => pgassign239,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign240,
      DIPB => net_gnd4,
      DOB => pgassign241,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign242
    );

  ramb16_30 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_30.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign243,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign244,
      DIPA => net_gnd4,
      DOA => pgassign245,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign246,
      ADDRB => pgassign247,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign248,
      DIPB => net_gnd4,
      DOB => pgassign249,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign250
    );

  ramb16_31 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_31.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign251,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign252,
      DIPA => net_gnd4,
      DOA => pgassign253,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign254,
      ADDRB => pgassign255,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign256,
      DIPB => net_gnd4,
      DOB => pgassign257,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign258
    );

  ramb16_32 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_32.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign259,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign260,
      DIPA => net_gnd4,
      DOA => pgassign261,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign262,
      ADDRB => pgassign263,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign264,
      DIPB => net_gnd4,
      DOB => pgassign265,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign266
    );

  ramb16_33 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_33.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign267,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign268,
      DIPA => net_gnd4,
      DOA => pgassign269,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign270,
      ADDRB => pgassign271,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign272,
      DIPB => net_gnd4,
      DOB => pgassign273,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign274
    );

  ramb16_34 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_34.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign275,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign276,
      DIPA => net_gnd4,
      DOA => pgassign277,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign278,
      ADDRB => pgassign279,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign280,
      DIPB => net_gnd4,
      DOB => pgassign281,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign282
    );

  ramb16_35 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_35.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign283,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign284,
      DIPA => net_gnd4,
      DOA => pgassign285,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign286,
      ADDRB => pgassign287,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign288,
      DIPB => net_gnd4,
      DOB => pgassign289,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign290
    );

  ramb16_36 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_36.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign291,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign292,
      DIPA => net_gnd4,
      DOA => pgassign293,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign294,
      ADDRB => pgassign295,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign296,
      DIPB => net_gnd4,
      DOB => pgassign297,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign298
    );

  ramb16_37 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_37.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign299,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign300,
      DIPA => net_gnd4,
      DOA => pgassign301,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign302,
      ADDRB => pgassign303,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign304,
      DIPB => net_gnd4,
      DOB => pgassign305,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign306
    );

  ramb16_38 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_38.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign307,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign308,
      DIPA => net_gnd4,
      DOA => pgassign309,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign310,
      ADDRB => pgassign311,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign312,
      DIPB => net_gnd4,
      DOB => pgassign313,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign314
    );

  ramb16_39 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_39.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign315,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign316,
      DIPA => net_gnd4,
      DOA => pgassign317,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign318,
      ADDRB => pgassign319,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign320,
      DIPB => net_gnd4,
      DOB => pgassign321,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign322
    );

  ramb16_40 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_40.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign323,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign324,
      DIPA => net_gnd4,
      DOA => pgassign325,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign326,
      ADDRB => pgassign327,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign328,
      DIPB => net_gnd4,
      DOB => pgassign329,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign330
    );

  ramb16_41 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_41.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign331,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign332,
      DIPA => net_gnd4,
      DOA => pgassign333,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign334,
      ADDRB => pgassign335,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign336,
      DIPB => net_gnd4,
      DOB => pgassign337,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign338
    );

  ramb16_42 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_42.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign339,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign340,
      DIPA => net_gnd4,
      DOA => pgassign341,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign342,
      ADDRB => pgassign343,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign344,
      DIPB => net_gnd4,
      DOB => pgassign345,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign346
    );

  ramb16_43 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_43.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign347,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign348,
      DIPA => net_gnd4,
      DOA => pgassign349,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign350,
      ADDRB => pgassign351,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign352,
      DIPB => net_gnd4,
      DOB => pgassign353,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign354
    );

  ramb16_44 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_44.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign355,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign356,
      DIPA => net_gnd4,
      DOA => pgassign357,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign358,
      ADDRB => pgassign359,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign360,
      DIPB => net_gnd4,
      DOB => pgassign361,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign362
    );

  ramb16_45 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_45.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign363,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign364,
      DIPA => net_gnd4,
      DOA => pgassign365,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign366,
      ADDRB => pgassign367,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign368,
      DIPB => net_gnd4,
      DOB => pgassign369,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign370
    );

  ramb16_46 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_46.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign371,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign372,
      DIPA => net_gnd4,
      DOA => pgassign373,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign374,
      ADDRB => pgassign375,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign376,
      DIPB => net_gnd4,
      DOB => pgassign377,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign378
    );

  ramb16_47 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_47.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign379,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign380,
      DIPA => net_gnd4,
      DOA => pgassign381,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign382,
      ADDRB => pgassign383,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign384,
      DIPB => net_gnd4,
      DOB => pgassign385,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign386
    );

  ramb16_48 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_48.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign387,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign388,
      DIPA => net_gnd4,
      DOA => pgassign389,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign390,
      ADDRB => pgassign391,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign392,
      DIPB => net_gnd4,
      DOB => pgassign393,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign394
    );

  ramb16_49 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_49.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign395,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign396,
      DIPA => net_gnd4,
      DOA => pgassign397,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign398,
      ADDRB => pgassign399,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign400,
      DIPB => net_gnd4,
      DOB => pgassign401,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign402
    );

  ramb16_50 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_50.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign403,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign404,
      DIPA => net_gnd4,
      DOA => pgassign405,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign406,
      ADDRB => pgassign407,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign408,
      DIPB => net_gnd4,
      DOB => pgassign409,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign410
    );

  ramb16_51 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_51.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign411,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign412,
      DIPA => net_gnd4,
      DOA => pgassign413,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign414,
      ADDRB => pgassign415,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign416,
      DIPB => net_gnd4,
      DOB => pgassign417,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign418
    );

  ramb16_52 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_52.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign419,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign420,
      DIPA => net_gnd4,
      DOA => pgassign421,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign422,
      ADDRB => pgassign423,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign424,
      DIPB => net_gnd4,
      DOB => pgassign425,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign426
    );

  ramb16_53 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_53.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign427,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign428,
      DIPA => net_gnd4,
      DOA => pgassign429,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign430,
      ADDRB => pgassign431,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign432,
      DIPB => net_gnd4,
      DOB => pgassign433,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign434
    );

  ramb16_54 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_54.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign435,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign436,
      DIPA => net_gnd4,
      DOA => pgassign437,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign438,
      ADDRB => pgassign439,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign440,
      DIPB => net_gnd4,
      DOB => pgassign441,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign442
    );

  ramb16_55 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_55.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign443,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign444,
      DIPA => net_gnd4,
      DOA => pgassign445,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign446,
      ADDRB => pgassign447,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign448,
      DIPB => net_gnd4,
      DOB => pgassign449,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign450
    );

  ramb16_56 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_56.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign451,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign452,
      DIPA => net_gnd4,
      DOA => pgassign453,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign454,
      ADDRB => pgassign455,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign456,
      DIPB => net_gnd4,
      DOB => pgassign457,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign458
    );

  ramb16_57 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_57.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign459,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign460,
      DIPA => net_gnd4,
      DOA => pgassign461,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign462,
      ADDRB => pgassign463,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign464,
      DIPB => net_gnd4,
      DOB => pgassign465,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign466
    );

  ramb16_58 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_58.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign467,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign468,
      DIPA => net_gnd4,
      DOA => pgassign469,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign470,
      ADDRB => pgassign471,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign472,
      DIPB => net_gnd4,
      DOB => pgassign473,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign474
    );

  ramb16_59 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_59.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign475,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign476,
      DIPA => net_gnd4,
      DOA => pgassign477,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign478,
      ADDRB => pgassign479,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign480,
      DIPB => net_gnd4,
      DOB => pgassign481,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign482
    );

  ramb16_60 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_60.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign483,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign484,
      DIPA => net_gnd4,
      DOA => pgassign485,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign486,
      ADDRB => pgassign487,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign488,
      DIPB => net_gnd4,
      DOB => pgassign489,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign490
    );

  ramb16_61 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_61.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign491,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign492,
      DIPA => net_gnd4,
      DOA => pgassign493,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign494,
      ADDRB => pgassign495,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign496,
      DIPB => net_gnd4,
      DOB => pgassign497,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign498
    );

  ramb16_62 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_62.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign499,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign500,
      DIPA => net_gnd4,
      DOA => pgassign501,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign502,
      ADDRB => pgassign503,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign504,
      DIPB => net_gnd4,
      DOB => pgassign505,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign506
    );

  ramb16_63 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_1_bram_combined_63.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign507,
      CASCADEINA => net_gnd0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign508,
      DIPA => net_gnd4,
      DOA => pgassign509,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign510,
      ADDRB => pgassign511,
      CASCADEINB => net_gnd0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign512,
      DIPB => net_gnd4,
      DOB => pgassign513,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign514
    );

end architecture STRUCTURE;

