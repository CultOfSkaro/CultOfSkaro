-------------------------------------------------------------------------------
-- plb_bram_if_cntlr_0_bram_elaborate.vhd
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

entity plb_bram_if_cntlr_0_bram_elaborate is
  generic (
    C_MEMSIZE : integer;
    C_PORT_DWIDTH : integer;
    C_PORT_AWIDTH : integer;
    C_NUM_WE : integer;
    C_FAMILY : string
    );
  port (
    BRAM_Rst_A : in std_logic;
    BRAM_Clk_A : in std_logic;
    BRAM_EN_A : in std_logic;
    BRAM_WEN_A : in std_logic_vector(0 to C_NUM_WE-1);
    BRAM_Addr_A : in std_logic_vector(0 to C_PORT_AWIDTH-1);
    BRAM_Din_A : out std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Dout_A : in std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Rst_B : in std_logic;
    BRAM_Clk_B : in std_logic;
    BRAM_EN_B : in std_logic;
    BRAM_WEN_B : in std_logic_vector(0 to C_NUM_WE-1);
    BRAM_Addr_B : in std_logic_vector(0 to C_PORT_AWIDTH-1);
    BRAM_Din_B : out std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Dout_B : in std_logic_vector(0 to C_PORT_DWIDTH-1)
  );

  attribute keep_hierarchy : STRING;
  attribute keep_hierarchy of plb_bram_if_cntlr_0_bram_elaborate : entity is "yes";

end plb_bram_if_cntlr_0_bram_elaborate;

architecture STRUCTURE of plb_bram_if_cntlr_0_bram_elaborate is

  component RAMB16 is
    generic (
      WRITE_MODE_A : string;
      WRITE_MODE_B : string;
      INIT_FILE : string;
      READ_WIDTH_A : integer;
      READ_WIDTH_B : integer;
      WRITE_WIDTH_A : integer;
      WRITE_WIDTH_B : integer;
      RAM_EXTENSION_A : string;
      RAM_EXTENSION_B : string
    );
    port (
      ADDRA : in std_logic_vector(14 downto 0);
      CASCADEINA : in std_logic;
      CASCADEOUTA : out std_logic;
      CLKA : in std_logic;
      DIA : in std_logic_vector(31 downto 0);
      DIPA : in std_logic_vector(3 downto 0);
      DOA : out std_logic_vector(31 downto 0);
      DOPA : out std_logic_vector(3 downto 0);
      ENA : in std_logic;
      REGCEA : in std_logic;
      SSRA : in std_logic;
      WEA : in std_logic_vector(3 downto 0);
      ADDRB : in std_logic_vector(14 downto 0);
      CASCADEINB : in std_logic;
      CASCADEOUTB : out std_logic;
      CLKB : in std_logic;
      DIB : in std_logic_vector(31 downto 0);
      DIPB : in std_logic_vector(3 downto 0);
      DOB : out std_logic_vector(31 downto 0);
      DOPB : out std_logic_vector(3 downto 0);
      ENB : in std_logic;
      REGCEB : in std_logic;
      SSRB : in std_logic;
      WEB : in std_logic_vector(3 downto 0)
    );
  end component;

  attribute BMM_INFO : STRING;

  attribute BMM_INFO of ramb16_0: label is " ";
  attribute BMM_INFO of ramb16_1: label is " ";
  attribute BMM_INFO of ramb16_2: label is " ";
  attribute BMM_INFO of ramb16_3: label is " ";
  attribute BMM_INFO of ramb16_4: label is " ";
  attribute BMM_INFO of ramb16_5: label is " ";
  attribute BMM_INFO of ramb16_6: label is " ";
  attribute BMM_INFO of ramb16_7: label is " ";
  attribute BMM_INFO of ramb16_8: label is " ";
  attribute BMM_INFO of ramb16_9: label is " ";
  attribute BMM_INFO of ramb16_10: label is " ";
  attribute BMM_INFO of ramb16_11: label is " ";
  attribute BMM_INFO of ramb16_12: label is " ";
  attribute BMM_INFO of ramb16_13: label is " ";
  attribute BMM_INFO of ramb16_14: label is " ";
  attribute BMM_INFO of ramb16_15: label is " ";
  attribute BMM_INFO of ramb16_16: label is " ";
  attribute BMM_INFO of ramb16_17: label is " ";
  attribute BMM_INFO of ramb16_18: label is " ";
  attribute BMM_INFO of ramb16_19: label is " ";
  attribute BMM_INFO of ramb16_20: label is " ";
  attribute BMM_INFO of ramb16_21: label is " ";
  attribute BMM_INFO of ramb16_22: label is " ";
  attribute BMM_INFO of ramb16_23: label is " ";
  attribute BMM_INFO of ramb16_24: label is " ";
  attribute BMM_INFO of ramb16_25: label is " ";
  attribute BMM_INFO of ramb16_26: label is " ";
  attribute BMM_INFO of ramb16_27: label is " ";
  attribute BMM_INFO of ramb16_28: label is " ";
  attribute BMM_INFO of ramb16_29: label is " ";
  attribute BMM_INFO of ramb16_30: label is " ";
  attribute BMM_INFO of ramb16_31: label is " ";
  attribute BMM_INFO of ramb16_32: label is " ";
  attribute BMM_INFO of ramb16_33: label is " ";
  attribute BMM_INFO of ramb16_34: label is " ";
  attribute BMM_INFO of ramb16_35: label is " ";
  attribute BMM_INFO of ramb16_36: label is " ";
  attribute BMM_INFO of ramb16_37: label is " ";
  attribute BMM_INFO of ramb16_38: label is " ";
  attribute BMM_INFO of ramb16_39: label is " ";
  attribute BMM_INFO of ramb16_40: label is " ";
  attribute BMM_INFO of ramb16_41: label is " ";
  attribute BMM_INFO of ramb16_42: label is " ";
  attribute BMM_INFO of ramb16_43: label is " ";
  attribute BMM_INFO of ramb16_44: label is " ";
  attribute BMM_INFO of ramb16_45: label is " ";
  attribute BMM_INFO of ramb16_46: label is " ";
  attribute BMM_INFO of ramb16_47: label is " ";
  attribute BMM_INFO of ramb16_48: label is " ";
  attribute BMM_INFO of ramb16_49: label is " ";
  attribute BMM_INFO of ramb16_50: label is " ";
  attribute BMM_INFO of ramb16_51: label is " ";
  attribute BMM_INFO of ramb16_52: label is " ";
  attribute BMM_INFO of ramb16_53: label is " ";
  attribute BMM_INFO of ramb16_54: label is " ";
  attribute BMM_INFO of ramb16_55: label is " ";
  attribute BMM_INFO of ramb16_56: label is " ";
  attribute BMM_INFO of ramb16_57: label is " ";
  attribute BMM_INFO of ramb16_58: label is " ";
  attribute BMM_INFO of ramb16_59: label is " ";
  attribute BMM_INFO of ramb16_60: label is " ";
  attribute BMM_INFO of ramb16_61: label is " ";
  attribute BMM_INFO of ramb16_62: label is " ";
  attribute BMM_INFO of ramb16_63: label is " ";
  attribute BMM_INFO of ramb16_64: label is " ";
  attribute BMM_INFO of ramb16_65: label is " ";
  attribute BMM_INFO of ramb16_66: label is " ";
  attribute BMM_INFO of ramb16_67: label is " ";
  attribute BMM_INFO of ramb16_68: label is " ";
  attribute BMM_INFO of ramb16_69: label is " ";
  attribute BMM_INFO of ramb16_70: label is " ";
  attribute BMM_INFO of ramb16_71: label is " ";
  attribute BMM_INFO of ramb16_72: label is " ";
  attribute BMM_INFO of ramb16_73: label is " ";
  attribute BMM_INFO of ramb16_74: label is " ";
  attribute BMM_INFO of ramb16_75: label is " ";
  attribute BMM_INFO of ramb16_76: label is " ";
  attribute BMM_INFO of ramb16_77: label is " ";
  attribute BMM_INFO of ramb16_78: label is " ";
  attribute BMM_INFO of ramb16_79: label is " ";
  attribute BMM_INFO of ramb16_80: label is " ";
  attribute BMM_INFO of ramb16_81: label is " ";
  attribute BMM_INFO of ramb16_82: label is " ";
  attribute BMM_INFO of ramb16_83: label is " ";
  attribute BMM_INFO of ramb16_84: label is " ";
  attribute BMM_INFO of ramb16_85: label is " ";
  attribute BMM_INFO of ramb16_86: label is " ";
  attribute BMM_INFO of ramb16_87: label is " ";
  attribute BMM_INFO of ramb16_88: label is " ";
  attribute BMM_INFO of ramb16_89: label is " ";
  attribute BMM_INFO of ramb16_90: label is " ";
  attribute BMM_INFO of ramb16_91: label is " ";
  attribute BMM_INFO of ramb16_92: label is " ";
  attribute BMM_INFO of ramb16_93: label is " ";
  attribute BMM_INFO of ramb16_94: label is " ";
  attribute BMM_INFO of ramb16_95: label is " ";
  attribute BMM_INFO of ramb16_96: label is " ";
  attribute BMM_INFO of ramb16_97: label is " ";
  attribute BMM_INFO of ramb16_98: label is " ";
  attribute BMM_INFO of ramb16_99: label is " ";
  attribute BMM_INFO of ramb16_100: label is " ";
  attribute BMM_INFO of ramb16_101: label is " ";
  attribute BMM_INFO of ramb16_102: label is " ";
  attribute BMM_INFO of ramb16_103: label is " ";
  attribute BMM_INFO of ramb16_104: label is " ";
  attribute BMM_INFO of ramb16_105: label is " ";
  attribute BMM_INFO of ramb16_106: label is " ";
  attribute BMM_INFO of ramb16_107: label is " ";
  attribute BMM_INFO of ramb16_108: label is " ";
  attribute BMM_INFO of ramb16_109: label is " ";
  attribute BMM_INFO of ramb16_110: label is " ";
  attribute BMM_INFO of ramb16_111: label is " ";
  attribute BMM_INFO of ramb16_112: label is " ";
  attribute BMM_INFO of ramb16_113: label is " ";
  attribute BMM_INFO of ramb16_114: label is " ";
  attribute BMM_INFO of ramb16_115: label is " ";
  attribute BMM_INFO of ramb16_116: label is " ";
  attribute BMM_INFO of ramb16_117: label is " ";
  attribute BMM_INFO of ramb16_118: label is " ";
  attribute BMM_INFO of ramb16_119: label is " ";
  attribute BMM_INFO of ramb16_120: label is " ";
  attribute BMM_INFO of ramb16_121: label is " ";
  attribute BMM_INFO of ramb16_122: label is " ";
  attribute BMM_INFO of ramb16_123: label is " ";
  attribute BMM_INFO of ramb16_124: label is " ";
  attribute BMM_INFO of ramb16_125: label is " ";
  attribute BMM_INFO of ramb16_126: label is " ";
  attribute BMM_INFO of ramb16_127: label is " ";
  -- Internal signals

  signal CASCADEA_0 : std_logic;
  signal CASCADEA_1 : std_logic;
  signal CASCADEA_2 : std_logic;
  signal CASCADEA_3 : std_logic;
  signal CASCADEA_4 : std_logic;
  signal CASCADEA_5 : std_logic;
  signal CASCADEA_6 : std_logic;
  signal CASCADEA_7 : std_logic;
  signal CASCADEA_8 : std_logic;
  signal CASCADEA_9 : std_logic;
  signal CASCADEA_10 : std_logic;
  signal CASCADEA_11 : std_logic;
  signal CASCADEA_12 : std_logic;
  signal CASCADEA_13 : std_logic;
  signal CASCADEA_14 : std_logic;
  signal CASCADEA_15 : std_logic;
  signal CASCADEA_16 : std_logic;
  signal CASCADEA_17 : std_logic;
  signal CASCADEA_18 : std_logic;
  signal CASCADEA_19 : std_logic;
  signal CASCADEA_20 : std_logic;
  signal CASCADEA_21 : std_logic;
  signal CASCADEA_22 : std_logic;
  signal CASCADEA_23 : std_logic;
  signal CASCADEA_24 : std_logic;
  signal CASCADEA_25 : std_logic;
  signal CASCADEA_26 : std_logic;
  signal CASCADEA_27 : std_logic;
  signal CASCADEA_28 : std_logic;
  signal CASCADEA_29 : std_logic;
  signal CASCADEA_30 : std_logic;
  signal CASCADEA_31 : std_logic;
  signal CASCADEA_32 : std_logic;
  signal CASCADEA_33 : std_logic;
  signal CASCADEA_34 : std_logic;
  signal CASCADEA_35 : std_logic;
  signal CASCADEA_36 : std_logic;
  signal CASCADEA_37 : std_logic;
  signal CASCADEA_38 : std_logic;
  signal CASCADEA_39 : std_logic;
  signal CASCADEA_40 : std_logic;
  signal CASCADEA_41 : std_logic;
  signal CASCADEA_42 : std_logic;
  signal CASCADEA_43 : std_logic;
  signal CASCADEA_44 : std_logic;
  signal CASCADEA_45 : std_logic;
  signal CASCADEA_46 : std_logic;
  signal CASCADEA_47 : std_logic;
  signal CASCADEA_48 : std_logic;
  signal CASCADEA_49 : std_logic;
  signal CASCADEA_50 : std_logic;
  signal CASCADEA_51 : std_logic;
  signal CASCADEA_52 : std_logic;
  signal CASCADEA_53 : std_logic;
  signal CASCADEA_54 : std_logic;
  signal CASCADEA_55 : std_logic;
  signal CASCADEA_56 : std_logic;
  signal CASCADEA_57 : std_logic;
  signal CASCADEA_58 : std_logic;
  signal CASCADEA_59 : std_logic;
  signal CASCADEA_60 : std_logic;
  signal CASCADEA_61 : std_logic;
  signal CASCADEA_62 : std_logic;
  signal CASCADEA_63 : std_logic;
  signal CASCADEB_0 : std_logic;
  signal CASCADEB_1 : std_logic;
  signal CASCADEB_2 : std_logic;
  signal CASCADEB_3 : std_logic;
  signal CASCADEB_4 : std_logic;
  signal CASCADEB_5 : std_logic;
  signal CASCADEB_6 : std_logic;
  signal CASCADEB_7 : std_logic;
  signal CASCADEB_8 : std_logic;
  signal CASCADEB_9 : std_logic;
  signal CASCADEB_10 : std_logic;
  signal CASCADEB_11 : std_logic;
  signal CASCADEB_12 : std_logic;
  signal CASCADEB_13 : std_logic;
  signal CASCADEB_14 : std_logic;
  signal CASCADEB_15 : std_logic;
  signal CASCADEB_16 : std_logic;
  signal CASCADEB_17 : std_logic;
  signal CASCADEB_18 : std_logic;
  signal CASCADEB_19 : std_logic;
  signal CASCADEB_20 : std_logic;
  signal CASCADEB_21 : std_logic;
  signal CASCADEB_22 : std_logic;
  signal CASCADEB_23 : std_logic;
  signal CASCADEB_24 : std_logic;
  signal CASCADEB_25 : std_logic;
  signal CASCADEB_26 : std_logic;
  signal CASCADEB_27 : std_logic;
  signal CASCADEB_28 : std_logic;
  signal CASCADEB_29 : std_logic;
  signal CASCADEB_30 : std_logic;
  signal CASCADEB_31 : std_logic;
  signal CASCADEB_32 : std_logic;
  signal CASCADEB_33 : std_logic;
  signal CASCADEB_34 : std_logic;
  signal CASCADEB_35 : std_logic;
  signal CASCADEB_36 : std_logic;
  signal CASCADEB_37 : std_logic;
  signal CASCADEB_38 : std_logic;
  signal CASCADEB_39 : std_logic;
  signal CASCADEB_40 : std_logic;
  signal CASCADEB_41 : std_logic;
  signal CASCADEB_42 : std_logic;
  signal CASCADEB_43 : std_logic;
  signal CASCADEB_44 : std_logic;
  signal CASCADEB_45 : std_logic;
  signal CASCADEB_46 : std_logic;
  signal CASCADEB_47 : std_logic;
  signal CASCADEB_48 : std_logic;
  signal CASCADEB_49 : std_logic;
  signal CASCADEB_50 : std_logic;
  signal CASCADEB_51 : std_logic;
  signal CASCADEB_52 : std_logic;
  signal CASCADEB_53 : std_logic;
  signal CASCADEB_54 : std_logic;
  signal CASCADEB_55 : std_logic;
  signal CASCADEB_56 : std_logic;
  signal CASCADEB_57 : std_logic;
  signal CASCADEB_58 : std_logic;
  signal CASCADEB_59 : std_logic;
  signal CASCADEB_60 : std_logic;
  signal CASCADEB_61 : std_logic;
  signal CASCADEB_62 : std_logic;
  signal CASCADEB_63 : std_logic;
  signal net_gnd0 : std_logic;
  signal net_gnd4 : std_logic_vector(3 downto 0);
  signal pgassign1 : std_logic_vector(0 to 30);
  signal pgassign2 : std_logic_vector(31 downto 0);
  signal pgassign3 : std_logic_vector(3 downto 0);
  signal pgassign4 : std_logic_vector(31 downto 0);
  signal pgassign5 : std_logic_vector(3 downto 0);
  signal pgassign6 : std_logic_vector(31 downto 0);
  signal pgassign7 : std_logic_vector(3 downto 0);
  signal pgassign8 : std_logic_vector(31 downto 0);
  signal pgassign9 : std_logic_vector(3 downto 0);
  signal pgassign10 : std_logic_vector(31 downto 0);
  signal pgassign11 : std_logic_vector(3 downto 0);
  signal pgassign12 : std_logic_vector(31 downto 0);
  signal pgassign13 : std_logic_vector(3 downto 0);
  signal pgassign14 : std_logic_vector(31 downto 0);
  signal pgassign15 : std_logic_vector(3 downto 0);
  signal pgassign16 : std_logic_vector(31 downto 0);
  signal pgassign17 : std_logic_vector(3 downto 0);
  signal pgassign18 : std_logic_vector(31 downto 0);
  signal pgassign19 : std_logic_vector(3 downto 0);
  signal pgassign20 : std_logic_vector(31 downto 0);
  signal pgassign21 : std_logic_vector(3 downto 0);
  signal pgassign22 : std_logic_vector(31 downto 0);
  signal pgassign23 : std_logic_vector(3 downto 0);
  signal pgassign24 : std_logic_vector(31 downto 0);
  signal pgassign25 : std_logic_vector(3 downto 0);
  signal pgassign26 : std_logic_vector(31 downto 0);
  signal pgassign27 : std_logic_vector(3 downto 0);
  signal pgassign28 : std_logic_vector(31 downto 0);
  signal pgassign29 : std_logic_vector(3 downto 0);
  signal pgassign30 : std_logic_vector(31 downto 0);
  signal pgassign31 : std_logic_vector(3 downto 0);
  signal pgassign32 : std_logic_vector(31 downto 0);
  signal pgassign33 : std_logic_vector(3 downto 0);
  signal pgassign34 : std_logic_vector(31 downto 0);
  signal pgassign35 : std_logic_vector(3 downto 0);
  signal pgassign36 : std_logic_vector(31 downto 0);
  signal pgassign37 : std_logic_vector(3 downto 0);
  signal pgassign38 : std_logic_vector(31 downto 0);
  signal pgassign39 : std_logic_vector(3 downto 0);
  signal pgassign40 : std_logic_vector(31 downto 0);
  signal pgassign41 : std_logic_vector(3 downto 0);
  signal pgassign42 : std_logic_vector(31 downto 0);
  signal pgassign43 : std_logic_vector(3 downto 0);
  signal pgassign44 : std_logic_vector(31 downto 0);
  signal pgassign45 : std_logic_vector(3 downto 0);
  signal pgassign46 : std_logic_vector(31 downto 0);
  signal pgassign47 : std_logic_vector(3 downto 0);
  signal pgassign48 : std_logic_vector(31 downto 0);
  signal pgassign49 : std_logic_vector(3 downto 0);
  signal pgassign50 : std_logic_vector(31 downto 0);
  signal pgassign51 : std_logic_vector(3 downto 0);
  signal pgassign52 : std_logic_vector(31 downto 0);
  signal pgassign53 : std_logic_vector(3 downto 0);
  signal pgassign54 : std_logic_vector(31 downto 0);
  signal pgassign55 : std_logic_vector(3 downto 0);
  signal pgassign56 : std_logic_vector(31 downto 0);
  signal pgassign57 : std_logic_vector(3 downto 0);
  signal pgassign58 : std_logic_vector(31 downto 0);
  signal pgassign59 : std_logic_vector(3 downto 0);
  signal pgassign60 : std_logic_vector(31 downto 0);
  signal pgassign61 : std_logic_vector(3 downto 0);
  signal pgassign62 : std_logic_vector(31 downto 0);
  signal pgassign63 : std_logic_vector(3 downto 0);
  signal pgassign64 : std_logic_vector(31 downto 0);
  signal pgassign65 : std_logic_vector(3 downto 0);
  signal pgassign66 : std_logic_vector(31 downto 0);
  signal pgassign67 : std_logic_vector(3 downto 0);
  signal pgassign68 : std_logic_vector(31 downto 0);
  signal pgassign69 : std_logic_vector(3 downto 0);
  signal pgassign70 : std_logic_vector(31 downto 0);
  signal pgassign71 : std_logic_vector(3 downto 0);
  signal pgassign72 : std_logic_vector(31 downto 0);
  signal pgassign73 : std_logic_vector(3 downto 0);
  signal pgassign74 : std_logic_vector(31 downto 0);
  signal pgassign75 : std_logic_vector(3 downto 0);
  signal pgassign76 : std_logic_vector(31 downto 0);
  signal pgassign77 : std_logic_vector(3 downto 0);
  signal pgassign78 : std_logic_vector(31 downto 0);
  signal pgassign79 : std_logic_vector(3 downto 0);
  signal pgassign80 : std_logic_vector(31 downto 0);
  signal pgassign81 : std_logic_vector(3 downto 0);
  signal pgassign82 : std_logic_vector(31 downto 0);
  signal pgassign83 : std_logic_vector(3 downto 0);
  signal pgassign84 : std_logic_vector(31 downto 0);
  signal pgassign85 : std_logic_vector(3 downto 0);
  signal pgassign86 : std_logic_vector(31 downto 0);
  signal pgassign87 : std_logic_vector(3 downto 0);
  signal pgassign88 : std_logic_vector(31 downto 0);
  signal pgassign89 : std_logic_vector(3 downto 0);
  signal pgassign90 : std_logic_vector(31 downto 0);
  signal pgassign91 : std_logic_vector(3 downto 0);
  signal pgassign92 : std_logic_vector(31 downto 0);
  signal pgassign93 : std_logic_vector(3 downto 0);
  signal pgassign94 : std_logic_vector(31 downto 0);
  signal pgassign95 : std_logic_vector(3 downto 0);
  signal pgassign96 : std_logic_vector(31 downto 0);
  signal pgassign97 : std_logic_vector(3 downto 0);
  signal pgassign98 : std_logic_vector(31 downto 0);
  signal pgassign99 : std_logic_vector(3 downto 0);
  signal pgassign100 : std_logic_vector(31 downto 0);
  signal pgassign101 : std_logic_vector(3 downto 0);
  signal pgassign102 : std_logic_vector(31 downto 0);
  signal pgassign103 : std_logic_vector(3 downto 0);
  signal pgassign104 : std_logic_vector(31 downto 0);
  signal pgassign105 : std_logic_vector(3 downto 0);
  signal pgassign106 : std_logic_vector(31 downto 0);
  signal pgassign107 : std_logic_vector(3 downto 0);
  signal pgassign108 : std_logic_vector(31 downto 0);
  signal pgassign109 : std_logic_vector(3 downto 0);
  signal pgassign110 : std_logic_vector(31 downto 0);
  signal pgassign111 : std_logic_vector(3 downto 0);
  signal pgassign112 : std_logic_vector(31 downto 0);
  signal pgassign113 : std_logic_vector(3 downto 0);
  signal pgassign114 : std_logic_vector(31 downto 0);
  signal pgassign115 : std_logic_vector(3 downto 0);
  signal pgassign116 : std_logic_vector(31 downto 0);
  signal pgassign117 : std_logic_vector(3 downto 0);
  signal pgassign118 : std_logic_vector(31 downto 0);
  signal pgassign119 : std_logic_vector(3 downto 0);
  signal pgassign120 : std_logic_vector(31 downto 0);
  signal pgassign121 : std_logic_vector(3 downto 0);
  signal pgassign122 : std_logic_vector(31 downto 0);
  signal pgassign123 : std_logic_vector(3 downto 0);
  signal pgassign124 : std_logic_vector(31 downto 0);
  signal pgassign125 : std_logic_vector(3 downto 0);
  signal pgassign126 : std_logic_vector(31 downto 0);
  signal pgassign127 : std_logic_vector(3 downto 0);
  signal pgassign128 : std_logic_vector(31 downto 0);
  signal pgassign129 : std_logic_vector(3 downto 0);
  signal pgassign130 : std_logic_vector(31 downto 0);
  signal pgassign131 : std_logic_vector(3 downto 0);
  signal pgassign132 : std_logic_vector(31 downto 0);
  signal pgassign133 : std_logic_vector(3 downto 0);
  signal pgassign134 : std_logic_vector(31 downto 0);
  signal pgassign135 : std_logic_vector(3 downto 0);
  signal pgassign136 : std_logic_vector(31 downto 0);
  signal pgassign137 : std_logic_vector(3 downto 0);
  signal pgassign138 : std_logic_vector(31 downto 0);
  signal pgassign139 : std_logic_vector(3 downto 0);
  signal pgassign140 : std_logic_vector(31 downto 0);
  signal pgassign141 : std_logic_vector(3 downto 0);
  signal pgassign142 : std_logic_vector(31 downto 0);
  signal pgassign143 : std_logic_vector(3 downto 0);
  signal pgassign144 : std_logic_vector(31 downto 0);
  signal pgassign145 : std_logic_vector(3 downto 0);
  signal pgassign146 : std_logic_vector(31 downto 0);
  signal pgassign147 : std_logic_vector(3 downto 0);
  signal pgassign148 : std_logic_vector(31 downto 0);
  signal pgassign149 : std_logic_vector(3 downto 0);
  signal pgassign150 : std_logic_vector(31 downto 0);
  signal pgassign151 : std_logic_vector(3 downto 0);
  signal pgassign152 : std_logic_vector(31 downto 0);
  signal pgassign153 : std_logic_vector(3 downto 0);
  signal pgassign154 : std_logic_vector(31 downto 0);
  signal pgassign155 : std_logic_vector(3 downto 0);
  signal pgassign156 : std_logic_vector(31 downto 0);
  signal pgassign157 : std_logic_vector(3 downto 0);
  signal pgassign158 : std_logic_vector(31 downto 0);
  signal pgassign159 : std_logic_vector(3 downto 0);
  signal pgassign160 : std_logic_vector(31 downto 0);
  signal pgassign161 : std_logic_vector(3 downto 0);
  signal pgassign162 : std_logic_vector(31 downto 0);
  signal pgassign163 : std_logic_vector(3 downto 0);
  signal pgassign164 : std_logic_vector(31 downto 0);
  signal pgassign165 : std_logic_vector(3 downto 0);
  signal pgassign166 : std_logic_vector(31 downto 0);
  signal pgassign167 : std_logic_vector(3 downto 0);
  signal pgassign168 : std_logic_vector(31 downto 0);
  signal pgassign169 : std_logic_vector(3 downto 0);
  signal pgassign170 : std_logic_vector(31 downto 0);
  signal pgassign171 : std_logic_vector(3 downto 0);
  signal pgassign172 : std_logic_vector(31 downto 0);
  signal pgassign173 : std_logic_vector(3 downto 0);
  signal pgassign174 : std_logic_vector(31 downto 0);
  signal pgassign175 : std_logic_vector(3 downto 0);
  signal pgassign176 : std_logic_vector(31 downto 0);
  signal pgassign177 : std_logic_vector(3 downto 0);
  signal pgassign178 : std_logic_vector(31 downto 0);
  signal pgassign179 : std_logic_vector(3 downto 0);
  signal pgassign180 : std_logic_vector(31 downto 0);
  signal pgassign181 : std_logic_vector(3 downto 0);
  signal pgassign182 : std_logic_vector(31 downto 0);
  signal pgassign183 : std_logic_vector(3 downto 0);
  signal pgassign184 : std_logic_vector(31 downto 0);
  signal pgassign185 : std_logic_vector(3 downto 0);
  signal pgassign186 : std_logic_vector(31 downto 0);
  signal pgassign187 : std_logic_vector(3 downto 0);
  signal pgassign188 : std_logic_vector(31 downto 0);
  signal pgassign189 : std_logic_vector(3 downto 0);
  signal pgassign190 : std_logic_vector(31 downto 0);
  signal pgassign191 : std_logic_vector(3 downto 0);
  signal pgassign192 : std_logic_vector(31 downto 0);
  signal pgassign193 : std_logic_vector(3 downto 0);
  signal pgassign194 : std_logic_vector(31 downto 0);
  signal pgassign195 : std_logic_vector(3 downto 0);
  signal pgassign196 : std_logic_vector(31 downto 0);
  signal pgassign197 : std_logic_vector(3 downto 0);
  signal pgassign198 : std_logic_vector(31 downto 0);
  signal pgassign199 : std_logic_vector(3 downto 0);
  signal pgassign200 : std_logic_vector(31 downto 0);
  signal pgassign201 : std_logic_vector(3 downto 0);
  signal pgassign202 : std_logic_vector(31 downto 0);
  signal pgassign203 : std_logic_vector(3 downto 0);
  signal pgassign204 : std_logic_vector(31 downto 0);
  signal pgassign205 : std_logic_vector(3 downto 0);
  signal pgassign206 : std_logic_vector(31 downto 0);
  signal pgassign207 : std_logic_vector(3 downto 0);
  signal pgassign208 : std_logic_vector(31 downto 0);
  signal pgassign209 : std_logic_vector(3 downto 0);
  signal pgassign210 : std_logic_vector(31 downto 0);
  signal pgassign211 : std_logic_vector(3 downto 0);
  signal pgassign212 : std_logic_vector(31 downto 0);
  signal pgassign213 : std_logic_vector(3 downto 0);
  signal pgassign214 : std_logic_vector(31 downto 0);
  signal pgassign215 : std_logic_vector(3 downto 0);
  signal pgassign216 : std_logic_vector(31 downto 0);
  signal pgassign217 : std_logic_vector(3 downto 0);
  signal pgassign218 : std_logic_vector(31 downto 0);
  signal pgassign219 : std_logic_vector(3 downto 0);
  signal pgassign220 : std_logic_vector(31 downto 0);
  signal pgassign221 : std_logic_vector(3 downto 0);
  signal pgassign222 : std_logic_vector(31 downto 0);
  signal pgassign223 : std_logic_vector(3 downto 0);
  signal pgassign224 : std_logic_vector(31 downto 0);
  signal pgassign225 : std_logic_vector(3 downto 0);
  signal pgassign226 : std_logic_vector(31 downto 0);
  signal pgassign227 : std_logic_vector(3 downto 0);
  signal pgassign228 : std_logic_vector(31 downto 0);
  signal pgassign229 : std_logic_vector(3 downto 0);
  signal pgassign230 : std_logic_vector(31 downto 0);
  signal pgassign231 : std_logic_vector(3 downto 0);
  signal pgassign232 : std_logic_vector(31 downto 0);
  signal pgassign233 : std_logic_vector(3 downto 0);
  signal pgassign234 : std_logic_vector(31 downto 0);
  signal pgassign235 : std_logic_vector(3 downto 0);
  signal pgassign236 : std_logic_vector(31 downto 0);
  signal pgassign237 : std_logic_vector(3 downto 0);
  signal pgassign238 : std_logic_vector(31 downto 0);
  signal pgassign239 : std_logic_vector(3 downto 0);
  signal pgassign240 : std_logic_vector(31 downto 0);
  signal pgassign241 : std_logic_vector(3 downto 0);
  signal pgassign242 : std_logic_vector(31 downto 0);
  signal pgassign243 : std_logic_vector(3 downto 0);
  signal pgassign244 : std_logic_vector(31 downto 0);
  signal pgassign245 : std_logic_vector(3 downto 0);
  signal pgassign246 : std_logic_vector(31 downto 0);
  signal pgassign247 : std_logic_vector(3 downto 0);
  signal pgassign248 : std_logic_vector(31 downto 0);
  signal pgassign249 : std_logic_vector(3 downto 0);
  signal pgassign250 : std_logic_vector(31 downto 0);
  signal pgassign251 : std_logic_vector(3 downto 0);
  signal pgassign252 : std_logic_vector(31 downto 0);
  signal pgassign253 : std_logic_vector(3 downto 0);
  signal pgassign254 : std_logic_vector(31 downto 0);
  signal pgassign255 : std_logic_vector(3 downto 0);
  signal pgassign256 : std_logic_vector(31 downto 0);
  signal pgassign257 : std_logic_vector(3 downto 0);
  signal pgassign258 : std_logic_vector(31 downto 0);
  signal pgassign259 : std_logic_vector(31 downto 0);
  signal pgassign260 : std_logic_vector(3 downto 0);
  signal pgassign261 : std_logic_vector(31 downto 0);
  signal pgassign262 : std_logic_vector(31 downto 0);
  signal pgassign263 : std_logic_vector(3 downto 0);
  signal pgassign264 : std_logic_vector(31 downto 0);
  signal pgassign265 : std_logic_vector(31 downto 0);
  signal pgassign266 : std_logic_vector(3 downto 0);
  signal pgassign267 : std_logic_vector(31 downto 0);
  signal pgassign268 : std_logic_vector(31 downto 0);
  signal pgassign269 : std_logic_vector(3 downto 0);
  signal pgassign270 : std_logic_vector(31 downto 0);
  signal pgassign271 : std_logic_vector(31 downto 0);
  signal pgassign272 : std_logic_vector(3 downto 0);
  signal pgassign273 : std_logic_vector(31 downto 0);
  signal pgassign274 : std_logic_vector(31 downto 0);
  signal pgassign275 : std_logic_vector(3 downto 0);
  signal pgassign276 : std_logic_vector(31 downto 0);
  signal pgassign277 : std_logic_vector(31 downto 0);
  signal pgassign278 : std_logic_vector(3 downto 0);
  signal pgassign279 : std_logic_vector(31 downto 0);
  signal pgassign280 : std_logic_vector(31 downto 0);
  signal pgassign281 : std_logic_vector(3 downto 0);
  signal pgassign282 : std_logic_vector(31 downto 0);
  signal pgassign283 : std_logic_vector(31 downto 0);
  signal pgassign284 : std_logic_vector(3 downto 0);
  signal pgassign285 : std_logic_vector(31 downto 0);
  signal pgassign286 : std_logic_vector(31 downto 0);
  signal pgassign287 : std_logic_vector(3 downto 0);
  signal pgassign288 : std_logic_vector(31 downto 0);
  signal pgassign289 : std_logic_vector(31 downto 0);
  signal pgassign290 : std_logic_vector(3 downto 0);
  signal pgassign291 : std_logic_vector(31 downto 0);
  signal pgassign292 : std_logic_vector(31 downto 0);
  signal pgassign293 : std_logic_vector(3 downto 0);
  signal pgassign294 : std_logic_vector(31 downto 0);
  signal pgassign295 : std_logic_vector(31 downto 0);
  signal pgassign296 : std_logic_vector(3 downto 0);
  signal pgassign297 : std_logic_vector(31 downto 0);
  signal pgassign298 : std_logic_vector(31 downto 0);
  signal pgassign299 : std_logic_vector(3 downto 0);
  signal pgassign300 : std_logic_vector(31 downto 0);
  signal pgassign301 : std_logic_vector(31 downto 0);
  signal pgassign302 : std_logic_vector(3 downto 0);
  signal pgassign303 : std_logic_vector(31 downto 0);
  signal pgassign304 : std_logic_vector(31 downto 0);
  signal pgassign305 : std_logic_vector(3 downto 0);
  signal pgassign306 : std_logic_vector(31 downto 0);
  signal pgassign307 : std_logic_vector(31 downto 0);
  signal pgassign308 : std_logic_vector(3 downto 0);
  signal pgassign309 : std_logic_vector(31 downto 0);
  signal pgassign310 : std_logic_vector(31 downto 0);
  signal pgassign311 : std_logic_vector(3 downto 0);
  signal pgassign312 : std_logic_vector(31 downto 0);
  signal pgassign313 : std_logic_vector(31 downto 0);
  signal pgassign314 : std_logic_vector(3 downto 0);
  signal pgassign315 : std_logic_vector(31 downto 0);
  signal pgassign316 : std_logic_vector(31 downto 0);
  signal pgassign317 : std_logic_vector(3 downto 0);
  signal pgassign318 : std_logic_vector(31 downto 0);
  signal pgassign319 : std_logic_vector(31 downto 0);
  signal pgassign320 : std_logic_vector(3 downto 0);
  signal pgassign321 : std_logic_vector(31 downto 0);
  signal pgassign322 : std_logic_vector(31 downto 0);
  signal pgassign323 : std_logic_vector(3 downto 0);
  signal pgassign324 : std_logic_vector(31 downto 0);
  signal pgassign325 : std_logic_vector(31 downto 0);
  signal pgassign326 : std_logic_vector(3 downto 0);
  signal pgassign327 : std_logic_vector(31 downto 0);
  signal pgassign328 : std_logic_vector(31 downto 0);
  signal pgassign329 : std_logic_vector(3 downto 0);
  signal pgassign330 : std_logic_vector(31 downto 0);
  signal pgassign331 : std_logic_vector(31 downto 0);
  signal pgassign332 : std_logic_vector(3 downto 0);
  signal pgassign333 : std_logic_vector(31 downto 0);
  signal pgassign334 : std_logic_vector(31 downto 0);
  signal pgassign335 : std_logic_vector(3 downto 0);
  signal pgassign336 : std_logic_vector(31 downto 0);
  signal pgassign337 : std_logic_vector(31 downto 0);
  signal pgassign338 : std_logic_vector(3 downto 0);
  signal pgassign339 : std_logic_vector(31 downto 0);
  signal pgassign340 : std_logic_vector(31 downto 0);
  signal pgassign341 : std_logic_vector(3 downto 0);
  signal pgassign342 : std_logic_vector(31 downto 0);
  signal pgassign343 : std_logic_vector(31 downto 0);
  signal pgassign344 : std_logic_vector(3 downto 0);
  signal pgassign345 : std_logic_vector(31 downto 0);
  signal pgassign346 : std_logic_vector(31 downto 0);
  signal pgassign347 : std_logic_vector(3 downto 0);
  signal pgassign348 : std_logic_vector(31 downto 0);
  signal pgassign349 : std_logic_vector(31 downto 0);
  signal pgassign350 : std_logic_vector(3 downto 0);
  signal pgassign351 : std_logic_vector(31 downto 0);
  signal pgassign352 : std_logic_vector(31 downto 0);
  signal pgassign353 : std_logic_vector(3 downto 0);
  signal pgassign354 : std_logic_vector(31 downto 0);
  signal pgassign355 : std_logic_vector(31 downto 0);
  signal pgassign356 : std_logic_vector(3 downto 0);
  signal pgassign357 : std_logic_vector(31 downto 0);
  signal pgassign358 : std_logic_vector(31 downto 0);
  signal pgassign359 : std_logic_vector(3 downto 0);
  signal pgassign360 : std_logic_vector(31 downto 0);
  signal pgassign361 : std_logic_vector(31 downto 0);
  signal pgassign362 : std_logic_vector(3 downto 0);
  signal pgassign363 : std_logic_vector(31 downto 0);
  signal pgassign364 : std_logic_vector(31 downto 0);
  signal pgassign365 : std_logic_vector(3 downto 0);
  signal pgassign366 : std_logic_vector(31 downto 0);
  signal pgassign367 : std_logic_vector(31 downto 0);
  signal pgassign368 : std_logic_vector(3 downto 0);
  signal pgassign369 : std_logic_vector(31 downto 0);
  signal pgassign370 : std_logic_vector(31 downto 0);
  signal pgassign371 : std_logic_vector(3 downto 0);
  signal pgassign372 : std_logic_vector(31 downto 0);
  signal pgassign373 : std_logic_vector(31 downto 0);
  signal pgassign374 : std_logic_vector(3 downto 0);
  signal pgassign375 : std_logic_vector(31 downto 0);
  signal pgassign376 : std_logic_vector(31 downto 0);
  signal pgassign377 : std_logic_vector(3 downto 0);
  signal pgassign378 : std_logic_vector(31 downto 0);
  signal pgassign379 : std_logic_vector(31 downto 0);
  signal pgassign380 : std_logic_vector(3 downto 0);
  signal pgassign381 : std_logic_vector(31 downto 0);
  signal pgassign382 : std_logic_vector(31 downto 0);
  signal pgassign383 : std_logic_vector(3 downto 0);
  signal pgassign384 : std_logic_vector(31 downto 0);
  signal pgassign385 : std_logic_vector(31 downto 0);
  signal pgassign386 : std_logic_vector(3 downto 0);
  signal pgassign387 : std_logic_vector(31 downto 0);
  signal pgassign388 : std_logic_vector(31 downto 0);
  signal pgassign389 : std_logic_vector(3 downto 0);
  signal pgassign390 : std_logic_vector(31 downto 0);
  signal pgassign391 : std_logic_vector(31 downto 0);
  signal pgassign392 : std_logic_vector(3 downto 0);
  signal pgassign393 : std_logic_vector(31 downto 0);
  signal pgassign394 : std_logic_vector(31 downto 0);
  signal pgassign395 : std_logic_vector(3 downto 0);
  signal pgassign396 : std_logic_vector(31 downto 0);
  signal pgassign397 : std_logic_vector(31 downto 0);
  signal pgassign398 : std_logic_vector(3 downto 0);
  signal pgassign399 : std_logic_vector(31 downto 0);
  signal pgassign400 : std_logic_vector(31 downto 0);
  signal pgassign401 : std_logic_vector(3 downto 0);
  signal pgassign402 : std_logic_vector(31 downto 0);
  signal pgassign403 : std_logic_vector(31 downto 0);
  signal pgassign404 : std_logic_vector(3 downto 0);
  signal pgassign405 : std_logic_vector(31 downto 0);
  signal pgassign406 : std_logic_vector(31 downto 0);
  signal pgassign407 : std_logic_vector(3 downto 0);
  signal pgassign408 : std_logic_vector(31 downto 0);
  signal pgassign409 : std_logic_vector(31 downto 0);
  signal pgassign410 : std_logic_vector(3 downto 0);
  signal pgassign411 : std_logic_vector(31 downto 0);
  signal pgassign412 : std_logic_vector(31 downto 0);
  signal pgassign413 : std_logic_vector(3 downto 0);
  signal pgassign414 : std_logic_vector(31 downto 0);
  signal pgassign415 : std_logic_vector(31 downto 0);
  signal pgassign416 : std_logic_vector(3 downto 0);
  signal pgassign417 : std_logic_vector(31 downto 0);
  signal pgassign418 : std_logic_vector(31 downto 0);
  signal pgassign419 : std_logic_vector(3 downto 0);
  signal pgassign420 : std_logic_vector(31 downto 0);
  signal pgassign421 : std_logic_vector(31 downto 0);
  signal pgassign422 : std_logic_vector(3 downto 0);
  signal pgassign423 : std_logic_vector(31 downto 0);
  signal pgassign424 : std_logic_vector(31 downto 0);
  signal pgassign425 : std_logic_vector(3 downto 0);
  signal pgassign426 : std_logic_vector(31 downto 0);
  signal pgassign427 : std_logic_vector(31 downto 0);
  signal pgassign428 : std_logic_vector(3 downto 0);
  signal pgassign429 : std_logic_vector(31 downto 0);
  signal pgassign430 : std_logic_vector(31 downto 0);
  signal pgassign431 : std_logic_vector(3 downto 0);
  signal pgassign432 : std_logic_vector(31 downto 0);
  signal pgassign433 : std_logic_vector(31 downto 0);
  signal pgassign434 : std_logic_vector(3 downto 0);
  signal pgassign435 : std_logic_vector(31 downto 0);
  signal pgassign436 : std_logic_vector(31 downto 0);
  signal pgassign437 : std_logic_vector(3 downto 0);
  signal pgassign438 : std_logic_vector(31 downto 0);
  signal pgassign439 : std_logic_vector(31 downto 0);
  signal pgassign440 : std_logic_vector(3 downto 0);
  signal pgassign441 : std_logic_vector(31 downto 0);
  signal pgassign442 : std_logic_vector(31 downto 0);
  signal pgassign443 : std_logic_vector(3 downto 0);
  signal pgassign444 : std_logic_vector(31 downto 0);
  signal pgassign445 : std_logic_vector(31 downto 0);
  signal pgassign446 : std_logic_vector(3 downto 0);
  signal pgassign447 : std_logic_vector(31 downto 0);
  signal pgassign448 : std_logic_vector(31 downto 0);
  signal pgassign449 : std_logic_vector(3 downto 0);
  signal pgassign450 : std_logic_vector(31 downto 0);
  signal pgassign451 : std_logic_vector(31 downto 0);
  signal pgassign452 : std_logic_vector(3 downto 0);
  signal pgassign453 : std_logic_vector(31 downto 0);
  signal pgassign454 : std_logic_vector(31 downto 0);
  signal pgassign455 : std_logic_vector(3 downto 0);
  signal pgassign456 : std_logic_vector(31 downto 0);
  signal pgassign457 : std_logic_vector(31 downto 0);
  signal pgassign458 : std_logic_vector(3 downto 0);
  signal pgassign459 : std_logic_vector(31 downto 0);
  signal pgassign460 : std_logic_vector(31 downto 0);
  signal pgassign461 : std_logic_vector(3 downto 0);
  signal pgassign462 : std_logic_vector(31 downto 0);
  signal pgassign463 : std_logic_vector(31 downto 0);
  signal pgassign464 : std_logic_vector(3 downto 0);
  signal pgassign465 : std_logic_vector(31 downto 0);
  signal pgassign466 : std_logic_vector(31 downto 0);
  signal pgassign467 : std_logic_vector(3 downto 0);
  signal pgassign468 : std_logic_vector(31 downto 0);
  signal pgassign469 : std_logic_vector(31 downto 0);
  signal pgassign470 : std_logic_vector(3 downto 0);
  signal pgassign471 : std_logic_vector(31 downto 0);
  signal pgassign472 : std_logic_vector(31 downto 0);
  signal pgassign473 : std_logic_vector(3 downto 0);
  signal pgassign474 : std_logic_vector(31 downto 0);
  signal pgassign475 : std_logic_vector(31 downto 0);
  signal pgassign476 : std_logic_vector(3 downto 0);
  signal pgassign477 : std_logic_vector(31 downto 0);
  signal pgassign478 : std_logic_vector(31 downto 0);
  signal pgassign479 : std_logic_vector(3 downto 0);
  signal pgassign480 : std_logic_vector(31 downto 0);
  signal pgassign481 : std_logic_vector(31 downto 0);
  signal pgassign482 : std_logic_vector(3 downto 0);
  signal pgassign483 : std_logic_vector(31 downto 0);
  signal pgassign484 : std_logic_vector(31 downto 0);
  signal pgassign485 : std_logic_vector(3 downto 0);
  signal pgassign486 : std_logic_vector(31 downto 0);
  signal pgassign487 : std_logic_vector(31 downto 0);
  signal pgassign488 : std_logic_vector(3 downto 0);
  signal pgassign489 : std_logic_vector(31 downto 0);
  signal pgassign490 : std_logic_vector(31 downto 0);
  signal pgassign491 : std_logic_vector(3 downto 0);
  signal pgassign492 : std_logic_vector(31 downto 0);
  signal pgassign493 : std_logic_vector(31 downto 0);
  signal pgassign494 : std_logic_vector(3 downto 0);
  signal pgassign495 : std_logic_vector(31 downto 0);
  signal pgassign496 : std_logic_vector(31 downto 0);
  signal pgassign497 : std_logic_vector(3 downto 0);
  signal pgassign498 : std_logic_vector(31 downto 0);
  signal pgassign499 : std_logic_vector(31 downto 0);
  signal pgassign500 : std_logic_vector(3 downto 0);
  signal pgassign501 : std_logic_vector(31 downto 0);
  signal pgassign502 : std_logic_vector(31 downto 0);
  signal pgassign503 : std_logic_vector(3 downto 0);
  signal pgassign504 : std_logic_vector(31 downto 0);
  signal pgassign505 : std_logic_vector(31 downto 0);
  signal pgassign506 : std_logic_vector(3 downto 0);
  signal pgassign507 : std_logic_vector(31 downto 0);
  signal pgassign508 : std_logic_vector(31 downto 0);
  signal pgassign509 : std_logic_vector(3 downto 0);
  signal pgassign510 : std_logic_vector(31 downto 0);
  signal pgassign511 : std_logic_vector(31 downto 0);
  signal pgassign512 : std_logic_vector(3 downto 0);
  signal pgassign513 : std_logic_vector(31 downto 0);
  signal pgassign514 : std_logic_vector(31 downto 0);
  signal pgassign515 : std_logic_vector(3 downto 0);
  signal pgassign516 : std_logic_vector(31 downto 0);
  signal pgassign517 : std_logic_vector(31 downto 0);
  signal pgassign518 : std_logic_vector(3 downto 0);
  signal pgassign519 : std_logic_vector(31 downto 0);
  signal pgassign520 : std_logic_vector(31 downto 0);
  signal pgassign521 : std_logic_vector(3 downto 0);
  signal pgassign522 : std_logic_vector(31 downto 0);
  signal pgassign523 : std_logic_vector(31 downto 0);
  signal pgassign524 : std_logic_vector(3 downto 0);
  signal pgassign525 : std_logic_vector(31 downto 0);
  signal pgassign526 : std_logic_vector(31 downto 0);
  signal pgassign527 : std_logic_vector(3 downto 0);
  signal pgassign528 : std_logic_vector(31 downto 0);
  signal pgassign529 : std_logic_vector(31 downto 0);
  signal pgassign530 : std_logic_vector(3 downto 0);
  signal pgassign531 : std_logic_vector(31 downto 0);
  signal pgassign532 : std_logic_vector(31 downto 0);
  signal pgassign533 : std_logic_vector(3 downto 0);
  signal pgassign534 : std_logic_vector(31 downto 0);
  signal pgassign535 : std_logic_vector(31 downto 0);
  signal pgassign536 : std_logic_vector(3 downto 0);
  signal pgassign537 : std_logic_vector(31 downto 0);
  signal pgassign538 : std_logic_vector(31 downto 0);
  signal pgassign539 : std_logic_vector(3 downto 0);
  signal pgassign540 : std_logic_vector(31 downto 0);
  signal pgassign541 : std_logic_vector(31 downto 0);
  signal pgassign542 : std_logic_vector(3 downto 0);
  signal pgassign543 : std_logic_vector(31 downto 0);
  signal pgassign544 : std_logic_vector(31 downto 0);
  signal pgassign545 : std_logic_vector(3 downto 0);
  signal pgassign546 : std_logic_vector(31 downto 0);
  signal pgassign547 : std_logic_vector(31 downto 0);
  signal pgassign548 : std_logic_vector(3 downto 0);
  signal pgassign549 : std_logic_vector(31 downto 0);
  signal pgassign550 : std_logic_vector(31 downto 0);
  signal pgassign551 : std_logic_vector(3 downto 0);
  signal pgassign552 : std_logic_vector(31 downto 0);
  signal pgassign553 : std_logic_vector(31 downto 0);
  signal pgassign554 : std_logic_vector(3 downto 0);
  signal pgassign555 : std_logic_vector(31 downto 0);
  signal pgassign556 : std_logic_vector(31 downto 0);
  signal pgassign557 : std_logic_vector(3 downto 0);
  signal pgassign558 : std_logic_vector(31 downto 0);
  signal pgassign559 : std_logic_vector(31 downto 0);
  signal pgassign560 : std_logic_vector(3 downto 0);
  signal pgassign561 : std_logic_vector(31 downto 0);
  signal pgassign562 : std_logic_vector(31 downto 0);
  signal pgassign563 : std_logic_vector(3 downto 0);
  signal pgassign564 : std_logic_vector(31 downto 0);
  signal pgassign565 : std_logic_vector(31 downto 0);
  signal pgassign566 : std_logic_vector(3 downto 0);
  signal pgassign567 : std_logic_vector(31 downto 0);
  signal pgassign568 : std_logic_vector(31 downto 0);
  signal pgassign569 : std_logic_vector(3 downto 0);
  signal pgassign570 : std_logic_vector(31 downto 0);
  signal pgassign571 : std_logic_vector(31 downto 0);
  signal pgassign572 : std_logic_vector(3 downto 0);
  signal pgassign573 : std_logic_vector(31 downto 0);
  signal pgassign574 : std_logic_vector(31 downto 0);
  signal pgassign575 : std_logic_vector(3 downto 0);
  signal pgassign576 : std_logic_vector(31 downto 0);
  signal pgassign577 : std_logic_vector(31 downto 0);
  signal pgassign578 : std_logic_vector(3 downto 0);
  signal pgassign579 : std_logic_vector(31 downto 0);
  signal pgassign580 : std_logic_vector(31 downto 0);
  signal pgassign581 : std_logic_vector(3 downto 0);
  signal pgassign582 : std_logic_vector(31 downto 0);
  signal pgassign583 : std_logic_vector(31 downto 0);
  signal pgassign584 : std_logic_vector(3 downto 0);
  signal pgassign585 : std_logic_vector(31 downto 0);
  signal pgassign586 : std_logic_vector(31 downto 0);
  signal pgassign587 : std_logic_vector(3 downto 0);
  signal pgassign588 : std_logic_vector(31 downto 0);
  signal pgassign589 : std_logic_vector(31 downto 0);
  signal pgassign590 : std_logic_vector(3 downto 0);
  signal pgassign591 : std_logic_vector(31 downto 0);
  signal pgassign592 : std_logic_vector(31 downto 0);
  signal pgassign593 : std_logic_vector(3 downto 0);
  signal pgassign594 : std_logic_vector(31 downto 0);
  signal pgassign595 : std_logic_vector(31 downto 0);
  signal pgassign596 : std_logic_vector(3 downto 0);
  signal pgassign597 : std_logic_vector(31 downto 0);
  signal pgassign598 : std_logic_vector(31 downto 0);
  signal pgassign599 : std_logic_vector(3 downto 0);
  signal pgassign600 : std_logic_vector(31 downto 0);
  signal pgassign601 : std_logic_vector(31 downto 0);
  signal pgassign602 : std_logic_vector(3 downto 0);
  signal pgassign603 : std_logic_vector(31 downto 0);
  signal pgassign604 : std_logic_vector(31 downto 0);
  signal pgassign605 : std_logic_vector(3 downto 0);
  signal pgassign606 : std_logic_vector(31 downto 0);
  signal pgassign607 : std_logic_vector(31 downto 0);
  signal pgassign608 : std_logic_vector(3 downto 0);
  signal pgassign609 : std_logic_vector(31 downto 0);
  signal pgassign610 : std_logic_vector(31 downto 0);
  signal pgassign611 : std_logic_vector(3 downto 0);
  signal pgassign612 : std_logic_vector(31 downto 0);
  signal pgassign613 : std_logic_vector(31 downto 0);
  signal pgassign614 : std_logic_vector(3 downto 0);
  signal pgassign615 : std_logic_vector(31 downto 0);
  signal pgassign616 : std_logic_vector(31 downto 0);
  signal pgassign617 : std_logic_vector(3 downto 0);
  signal pgassign618 : std_logic_vector(31 downto 0);
  signal pgassign619 : std_logic_vector(31 downto 0);
  signal pgassign620 : std_logic_vector(3 downto 0);
  signal pgassign621 : std_logic_vector(31 downto 0);
  signal pgassign622 : std_logic_vector(31 downto 0);
  signal pgassign623 : std_logic_vector(3 downto 0);
  signal pgassign624 : std_logic_vector(31 downto 0);
  signal pgassign625 : std_logic_vector(31 downto 0);
  signal pgassign626 : std_logic_vector(3 downto 0);
  signal pgassign627 : std_logic_vector(31 downto 0);
  signal pgassign628 : std_logic_vector(31 downto 0);
  signal pgassign629 : std_logic_vector(3 downto 0);
  signal pgassign630 : std_logic_vector(31 downto 0);
  signal pgassign631 : std_logic_vector(31 downto 0);
  signal pgassign632 : std_logic_vector(3 downto 0);
  signal pgassign633 : std_logic_vector(31 downto 0);
  signal pgassign634 : std_logic_vector(31 downto 0);
  signal pgassign635 : std_logic_vector(3 downto 0);
  signal pgassign636 : std_logic_vector(31 downto 0);
  signal pgassign637 : std_logic_vector(31 downto 0);
  signal pgassign638 : std_logic_vector(3 downto 0);
  signal pgassign639 : std_logic_vector(31 downto 0);
  signal pgassign640 : std_logic_vector(31 downto 0);
  signal pgassign641 : std_logic_vector(3 downto 0);

begin

  -- Internal assignments

  pgassign1(0 to 30) <= B"0000000000000000000000000000000";
  pgassign2(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign2(0 downto 0) <= BRAM_Dout_A(0 to 0);
  pgassign3(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign3(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign3(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign3(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign4(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign4(0 downto 0) <= BRAM_Dout_B(0 to 0);
  pgassign5(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign5(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign5(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign5(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign6(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign6(0 downto 0) <= BRAM_Dout_A(1 to 1);
  pgassign7(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign7(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign7(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign7(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign8(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign8(0 downto 0) <= BRAM_Dout_B(1 to 1);
  pgassign9(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign9(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign9(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign9(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign10(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign10(0 downto 0) <= BRAM_Dout_A(2 to 2);
  pgassign11(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign11(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign11(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign11(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign12(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign12(0 downto 0) <= BRAM_Dout_B(2 to 2);
  pgassign13(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign13(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign13(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign13(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign14(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign14(0 downto 0) <= BRAM_Dout_A(3 to 3);
  pgassign15(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign15(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign15(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign15(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign16(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign16(0 downto 0) <= BRAM_Dout_B(3 to 3);
  pgassign17(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign17(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign17(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign17(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign18(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign18(0 downto 0) <= BRAM_Dout_A(4 to 4);
  pgassign19(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign19(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign19(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign19(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign20(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign20(0 downto 0) <= BRAM_Dout_B(4 to 4);
  pgassign21(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign21(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign21(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign21(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign22(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign22(0 downto 0) <= BRAM_Dout_A(5 to 5);
  pgassign23(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign23(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign23(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign23(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign24(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign24(0 downto 0) <= BRAM_Dout_B(5 to 5);
  pgassign25(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign25(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign25(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign25(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign26(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign26(0 downto 0) <= BRAM_Dout_A(6 to 6);
  pgassign27(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign27(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign27(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign27(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign28(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign28(0 downto 0) <= BRAM_Dout_B(6 to 6);
  pgassign29(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign29(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign29(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign29(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign30(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign30(0 downto 0) <= BRAM_Dout_A(7 to 7);
  pgassign31(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign31(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign31(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign31(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign32(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign32(0 downto 0) <= BRAM_Dout_B(7 to 7);
  pgassign33(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign33(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign33(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign33(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign34(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign34(0 downto 0) <= BRAM_Dout_A(8 to 8);
  pgassign35(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign35(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign35(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign35(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign36(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign36(0 downto 0) <= BRAM_Dout_B(8 to 8);
  pgassign37(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign37(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign37(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign37(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign38(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign38(0 downto 0) <= BRAM_Dout_A(9 to 9);
  pgassign39(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign39(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign39(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign39(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign40(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign40(0 downto 0) <= BRAM_Dout_B(9 to 9);
  pgassign41(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign41(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign41(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign41(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign42(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign42(0 downto 0) <= BRAM_Dout_A(10 to 10);
  pgassign43(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign43(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign43(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign43(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign44(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign44(0 downto 0) <= BRAM_Dout_B(10 to 10);
  pgassign45(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign45(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign45(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign45(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign46(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign46(0 downto 0) <= BRAM_Dout_A(11 to 11);
  pgassign47(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign47(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign47(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign47(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign48(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign48(0 downto 0) <= BRAM_Dout_B(11 to 11);
  pgassign49(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign49(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign49(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign49(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign50(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign50(0 downto 0) <= BRAM_Dout_A(12 to 12);
  pgassign51(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign51(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign51(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign51(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign52(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign52(0 downto 0) <= BRAM_Dout_B(12 to 12);
  pgassign53(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign53(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign53(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign53(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign54(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign54(0 downto 0) <= BRAM_Dout_A(13 to 13);
  pgassign55(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign55(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign55(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign55(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign56(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign56(0 downto 0) <= BRAM_Dout_B(13 to 13);
  pgassign57(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign57(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign57(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign57(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign58(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign58(0 downto 0) <= BRAM_Dout_A(14 to 14);
  pgassign59(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign59(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign59(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign59(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign60(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign60(0 downto 0) <= BRAM_Dout_B(14 to 14);
  pgassign61(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign61(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign61(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign61(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign62(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign62(0 downto 0) <= BRAM_Dout_A(15 to 15);
  pgassign63(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign63(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign63(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign63(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign64(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign64(0 downto 0) <= BRAM_Dout_B(15 to 15);
  pgassign65(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign65(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign65(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign65(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign66(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign66(0 downto 0) <= BRAM_Dout_A(16 to 16);
  pgassign67(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign67(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign67(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign67(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign68(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign68(0 downto 0) <= BRAM_Dout_B(16 to 16);
  pgassign69(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign69(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign69(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign69(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign70(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign70(0 downto 0) <= BRAM_Dout_A(17 to 17);
  pgassign71(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign71(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign71(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign71(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign72(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign72(0 downto 0) <= BRAM_Dout_B(17 to 17);
  pgassign73(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign73(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign73(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign73(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign74(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign74(0 downto 0) <= BRAM_Dout_A(18 to 18);
  pgassign75(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign75(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign75(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign75(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign76(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign76(0 downto 0) <= BRAM_Dout_B(18 to 18);
  pgassign77(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign77(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign77(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign77(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign78(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign78(0 downto 0) <= BRAM_Dout_A(19 to 19);
  pgassign79(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign79(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign79(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign79(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign80(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign80(0 downto 0) <= BRAM_Dout_B(19 to 19);
  pgassign81(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign81(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign81(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign81(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign82(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign82(0 downto 0) <= BRAM_Dout_A(20 to 20);
  pgassign83(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign83(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign83(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign83(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign84(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign84(0 downto 0) <= BRAM_Dout_B(20 to 20);
  pgassign85(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign85(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign85(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign85(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign86(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign86(0 downto 0) <= BRAM_Dout_A(21 to 21);
  pgassign87(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign87(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign87(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign87(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign88(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign88(0 downto 0) <= BRAM_Dout_B(21 to 21);
  pgassign89(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign89(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign89(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign89(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign90(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign90(0 downto 0) <= BRAM_Dout_A(22 to 22);
  pgassign91(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign91(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign91(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign91(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign92(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign92(0 downto 0) <= BRAM_Dout_B(22 to 22);
  pgassign93(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign93(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign93(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign93(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign94(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign94(0 downto 0) <= BRAM_Dout_A(23 to 23);
  pgassign95(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign95(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign95(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign95(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign96(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign96(0 downto 0) <= BRAM_Dout_B(23 to 23);
  pgassign97(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign97(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign97(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign97(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign98(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign98(0 downto 0) <= BRAM_Dout_A(24 to 24);
  pgassign99(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign99(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign99(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign99(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign100(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign100(0 downto 0) <= BRAM_Dout_B(24 to 24);
  pgassign101(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign101(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign101(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign101(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign102(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign102(0 downto 0) <= BRAM_Dout_A(25 to 25);
  pgassign103(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign103(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign103(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign103(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign104(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign104(0 downto 0) <= BRAM_Dout_B(25 to 25);
  pgassign105(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign105(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign105(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign105(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign106(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign106(0 downto 0) <= BRAM_Dout_A(26 to 26);
  pgassign107(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign107(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign107(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign107(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign108(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign108(0 downto 0) <= BRAM_Dout_B(26 to 26);
  pgassign109(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign109(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign109(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign109(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign110(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign110(0 downto 0) <= BRAM_Dout_A(27 to 27);
  pgassign111(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign111(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign111(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign111(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign112(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign112(0 downto 0) <= BRAM_Dout_B(27 to 27);
  pgassign113(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign113(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign113(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign113(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign114(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign114(0 downto 0) <= BRAM_Dout_A(28 to 28);
  pgassign115(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign115(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign115(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign115(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign116(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign116(0 downto 0) <= BRAM_Dout_B(28 to 28);
  pgassign117(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign117(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign117(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign117(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign118(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign118(0 downto 0) <= BRAM_Dout_A(29 to 29);
  pgassign119(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign119(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign119(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign119(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign120(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign120(0 downto 0) <= BRAM_Dout_B(29 to 29);
  pgassign121(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign121(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign121(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign121(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign122(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign122(0 downto 0) <= BRAM_Dout_A(30 to 30);
  pgassign123(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign123(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign123(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign123(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign124(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign124(0 downto 0) <= BRAM_Dout_B(30 to 30);
  pgassign125(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign125(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign125(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign125(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign126(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign126(0 downto 0) <= BRAM_Dout_A(31 to 31);
  pgassign127(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign127(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign127(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign127(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign128(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign128(0 downto 0) <= BRAM_Dout_B(31 to 31);
  pgassign129(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign129(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign129(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign129(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign130(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign130(0 downto 0) <= BRAM_Dout_A(32 to 32);
  pgassign131(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign131(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign131(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign131(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign132(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign132(0 downto 0) <= BRAM_Dout_B(32 to 32);
  pgassign133(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign133(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign133(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign133(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign134(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign134(0 downto 0) <= BRAM_Dout_A(33 to 33);
  pgassign135(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign135(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign135(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign135(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign136(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign136(0 downto 0) <= BRAM_Dout_B(33 to 33);
  pgassign137(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign137(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign137(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign137(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign138(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign138(0 downto 0) <= BRAM_Dout_A(34 to 34);
  pgassign139(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign139(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign139(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign139(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign140(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign140(0 downto 0) <= BRAM_Dout_B(34 to 34);
  pgassign141(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign141(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign141(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign141(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign142(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign142(0 downto 0) <= BRAM_Dout_A(35 to 35);
  pgassign143(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign143(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign143(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign143(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign144(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign144(0 downto 0) <= BRAM_Dout_B(35 to 35);
  pgassign145(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign145(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign145(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign145(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign146(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign146(0 downto 0) <= BRAM_Dout_A(36 to 36);
  pgassign147(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign147(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign147(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign147(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign148(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign148(0 downto 0) <= BRAM_Dout_B(36 to 36);
  pgassign149(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign149(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign149(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign149(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign150(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign150(0 downto 0) <= BRAM_Dout_A(37 to 37);
  pgassign151(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign151(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign151(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign151(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign152(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign152(0 downto 0) <= BRAM_Dout_B(37 to 37);
  pgassign153(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign153(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign153(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign153(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign154(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign154(0 downto 0) <= BRAM_Dout_A(38 to 38);
  pgassign155(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign155(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign155(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign155(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign156(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign156(0 downto 0) <= BRAM_Dout_B(38 to 38);
  pgassign157(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign157(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign157(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign157(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign158(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign158(0 downto 0) <= BRAM_Dout_A(39 to 39);
  pgassign159(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign159(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign159(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign159(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign160(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign160(0 downto 0) <= BRAM_Dout_B(39 to 39);
  pgassign161(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign161(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign161(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign161(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign162(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign162(0 downto 0) <= BRAM_Dout_A(40 to 40);
  pgassign163(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign163(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign163(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign163(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign164(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign164(0 downto 0) <= BRAM_Dout_B(40 to 40);
  pgassign165(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign165(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign165(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign165(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign166(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign166(0 downto 0) <= BRAM_Dout_A(41 to 41);
  pgassign167(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign167(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign167(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign167(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign168(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign168(0 downto 0) <= BRAM_Dout_B(41 to 41);
  pgassign169(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign169(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign169(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign169(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign170(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign170(0 downto 0) <= BRAM_Dout_A(42 to 42);
  pgassign171(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign171(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign171(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign171(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign172(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign172(0 downto 0) <= BRAM_Dout_B(42 to 42);
  pgassign173(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign173(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign173(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign173(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign174(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign174(0 downto 0) <= BRAM_Dout_A(43 to 43);
  pgassign175(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign175(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign175(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign175(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign176(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign176(0 downto 0) <= BRAM_Dout_B(43 to 43);
  pgassign177(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign177(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign177(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign177(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign178(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign178(0 downto 0) <= BRAM_Dout_A(44 to 44);
  pgassign179(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign179(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign179(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign179(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign180(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign180(0 downto 0) <= BRAM_Dout_B(44 to 44);
  pgassign181(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign181(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign181(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign181(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign182(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign182(0 downto 0) <= BRAM_Dout_A(45 to 45);
  pgassign183(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign183(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign183(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign183(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign184(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign184(0 downto 0) <= BRAM_Dout_B(45 to 45);
  pgassign185(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign185(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign185(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign185(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign186(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign186(0 downto 0) <= BRAM_Dout_A(46 to 46);
  pgassign187(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign187(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign187(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign187(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign188(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign188(0 downto 0) <= BRAM_Dout_B(46 to 46);
  pgassign189(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign189(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign189(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign189(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign190(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign190(0 downto 0) <= BRAM_Dout_A(47 to 47);
  pgassign191(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign191(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign191(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign191(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign192(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign192(0 downto 0) <= BRAM_Dout_B(47 to 47);
  pgassign193(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign193(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign193(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign193(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign194(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign194(0 downto 0) <= BRAM_Dout_A(48 to 48);
  pgassign195(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign195(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign195(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign195(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign196(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign196(0 downto 0) <= BRAM_Dout_B(48 to 48);
  pgassign197(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign197(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign197(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign197(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign198(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign198(0 downto 0) <= BRAM_Dout_A(49 to 49);
  pgassign199(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign199(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign199(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign199(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign200(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign200(0 downto 0) <= BRAM_Dout_B(49 to 49);
  pgassign201(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign201(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign201(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign201(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign202(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign202(0 downto 0) <= BRAM_Dout_A(50 to 50);
  pgassign203(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign203(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign203(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign203(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign204(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign204(0 downto 0) <= BRAM_Dout_B(50 to 50);
  pgassign205(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign205(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign205(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign205(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign206(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign206(0 downto 0) <= BRAM_Dout_A(51 to 51);
  pgassign207(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign207(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign207(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign207(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign208(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign208(0 downto 0) <= BRAM_Dout_B(51 to 51);
  pgassign209(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign209(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign209(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign209(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign210(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign210(0 downto 0) <= BRAM_Dout_A(52 to 52);
  pgassign211(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign211(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign211(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign211(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign212(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign212(0 downto 0) <= BRAM_Dout_B(52 to 52);
  pgassign213(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign213(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign213(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign213(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign214(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign214(0 downto 0) <= BRAM_Dout_A(53 to 53);
  pgassign215(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign215(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign215(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign215(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign216(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign216(0 downto 0) <= BRAM_Dout_B(53 to 53);
  pgassign217(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign217(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign217(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign217(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign218(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign218(0 downto 0) <= BRAM_Dout_A(54 to 54);
  pgassign219(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign219(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign219(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign219(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign220(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign220(0 downto 0) <= BRAM_Dout_B(54 to 54);
  pgassign221(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign221(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign221(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign221(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign222(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign222(0 downto 0) <= BRAM_Dout_A(55 to 55);
  pgassign223(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign223(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign223(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign223(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign224(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign224(0 downto 0) <= BRAM_Dout_B(55 to 55);
  pgassign225(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign225(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign225(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign225(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign226(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign226(0 downto 0) <= BRAM_Dout_A(56 to 56);
  pgassign227(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign227(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign227(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign227(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign228(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign228(0 downto 0) <= BRAM_Dout_B(56 to 56);
  pgassign229(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign229(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign229(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign229(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign230(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign230(0 downto 0) <= BRAM_Dout_A(57 to 57);
  pgassign231(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign231(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign231(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign231(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign232(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign232(0 downto 0) <= BRAM_Dout_B(57 to 57);
  pgassign233(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign233(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign233(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign233(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign234(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign234(0 downto 0) <= BRAM_Dout_A(58 to 58);
  pgassign235(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign235(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign235(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign235(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign236(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign236(0 downto 0) <= BRAM_Dout_B(58 to 58);
  pgassign237(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign237(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign237(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign237(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign238(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign238(0 downto 0) <= BRAM_Dout_A(59 to 59);
  pgassign239(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign239(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign239(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign239(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign240(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign240(0 downto 0) <= BRAM_Dout_B(59 to 59);
  pgassign241(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign241(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign241(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign241(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign242(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign242(0 downto 0) <= BRAM_Dout_A(60 to 60);
  pgassign243(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign243(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign243(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign243(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign244(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign244(0 downto 0) <= BRAM_Dout_B(60 to 60);
  pgassign245(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign245(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign245(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign245(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign246(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign246(0 downto 0) <= BRAM_Dout_A(61 to 61);
  pgassign247(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign247(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign247(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign247(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign248(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign248(0 downto 0) <= BRAM_Dout_B(61 to 61);
  pgassign249(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign249(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign249(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign249(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign250(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign250(0 downto 0) <= BRAM_Dout_A(62 to 62);
  pgassign251(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign251(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign251(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign251(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign252(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign252(0 downto 0) <= BRAM_Dout_B(62 to 62);
  pgassign253(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign253(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign253(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign253(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign254(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign254(0 downto 0) <= BRAM_Dout_A(63 to 63);
  pgassign255(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign255(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign255(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign255(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign256(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign256(0 downto 0) <= BRAM_Dout_B(63 to 63);
  pgassign257(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign257(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign257(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign257(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign258(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign258(0 downto 0) <= BRAM_Dout_A(0 to 0);
  BRAM_Din_A(0 to 0) <= pgassign259(0 downto 0);
  pgassign260(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign260(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign260(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign260(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign261(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign261(0 downto 0) <= BRAM_Dout_B(0 to 0);
  BRAM_Din_B(0 to 0) <= pgassign262(0 downto 0);
  pgassign263(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign263(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign263(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign263(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign264(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign264(0 downto 0) <= BRAM_Dout_A(1 to 1);
  BRAM_Din_A(1 to 1) <= pgassign265(0 downto 0);
  pgassign266(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign266(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign266(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign266(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign267(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign267(0 downto 0) <= BRAM_Dout_B(1 to 1);
  BRAM_Din_B(1 to 1) <= pgassign268(0 downto 0);
  pgassign269(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign269(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign269(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign269(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign270(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign270(0 downto 0) <= BRAM_Dout_A(2 to 2);
  BRAM_Din_A(2 to 2) <= pgassign271(0 downto 0);
  pgassign272(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign272(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign272(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign272(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign273(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign273(0 downto 0) <= BRAM_Dout_B(2 to 2);
  BRAM_Din_B(2 to 2) <= pgassign274(0 downto 0);
  pgassign275(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign275(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign275(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign275(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign276(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign276(0 downto 0) <= BRAM_Dout_A(3 to 3);
  BRAM_Din_A(3 to 3) <= pgassign277(0 downto 0);
  pgassign278(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign278(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign278(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign278(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign279(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign279(0 downto 0) <= BRAM_Dout_B(3 to 3);
  BRAM_Din_B(3 to 3) <= pgassign280(0 downto 0);
  pgassign281(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign281(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign281(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign281(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign282(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign282(0 downto 0) <= BRAM_Dout_A(4 to 4);
  BRAM_Din_A(4 to 4) <= pgassign283(0 downto 0);
  pgassign284(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign284(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign284(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign284(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign285(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign285(0 downto 0) <= BRAM_Dout_B(4 to 4);
  BRAM_Din_B(4 to 4) <= pgassign286(0 downto 0);
  pgassign287(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign287(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign287(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign287(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign288(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign288(0 downto 0) <= BRAM_Dout_A(5 to 5);
  BRAM_Din_A(5 to 5) <= pgassign289(0 downto 0);
  pgassign290(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign290(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign290(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign290(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign291(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign291(0 downto 0) <= BRAM_Dout_B(5 to 5);
  BRAM_Din_B(5 to 5) <= pgassign292(0 downto 0);
  pgassign293(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign293(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign293(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign293(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign294(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign294(0 downto 0) <= BRAM_Dout_A(6 to 6);
  BRAM_Din_A(6 to 6) <= pgassign295(0 downto 0);
  pgassign296(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign296(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign296(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign296(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign297(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign297(0 downto 0) <= BRAM_Dout_B(6 to 6);
  BRAM_Din_B(6 to 6) <= pgassign298(0 downto 0);
  pgassign299(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign299(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign299(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign299(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign300(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign300(0 downto 0) <= BRAM_Dout_A(7 to 7);
  BRAM_Din_A(7 to 7) <= pgassign301(0 downto 0);
  pgassign302(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign302(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign302(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign302(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign303(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign303(0 downto 0) <= BRAM_Dout_B(7 to 7);
  BRAM_Din_B(7 to 7) <= pgassign304(0 downto 0);
  pgassign305(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign305(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign305(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign305(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign306(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign306(0 downto 0) <= BRAM_Dout_A(8 to 8);
  BRAM_Din_A(8 to 8) <= pgassign307(0 downto 0);
  pgassign308(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign308(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign308(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign308(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign309(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign309(0 downto 0) <= BRAM_Dout_B(8 to 8);
  BRAM_Din_B(8 to 8) <= pgassign310(0 downto 0);
  pgassign311(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign311(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign311(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign311(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign312(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign312(0 downto 0) <= BRAM_Dout_A(9 to 9);
  BRAM_Din_A(9 to 9) <= pgassign313(0 downto 0);
  pgassign314(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign314(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign314(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign314(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign315(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign315(0 downto 0) <= BRAM_Dout_B(9 to 9);
  BRAM_Din_B(9 to 9) <= pgassign316(0 downto 0);
  pgassign317(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign317(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign317(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign317(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign318(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign318(0 downto 0) <= BRAM_Dout_A(10 to 10);
  BRAM_Din_A(10 to 10) <= pgassign319(0 downto 0);
  pgassign320(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign320(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign320(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign320(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign321(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign321(0 downto 0) <= BRAM_Dout_B(10 to 10);
  BRAM_Din_B(10 to 10) <= pgassign322(0 downto 0);
  pgassign323(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign323(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign323(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign323(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign324(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign324(0 downto 0) <= BRAM_Dout_A(11 to 11);
  BRAM_Din_A(11 to 11) <= pgassign325(0 downto 0);
  pgassign326(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign326(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign326(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign326(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign327(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign327(0 downto 0) <= BRAM_Dout_B(11 to 11);
  BRAM_Din_B(11 to 11) <= pgassign328(0 downto 0);
  pgassign329(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign329(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign329(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign329(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign330(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign330(0 downto 0) <= BRAM_Dout_A(12 to 12);
  BRAM_Din_A(12 to 12) <= pgassign331(0 downto 0);
  pgassign332(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign332(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign332(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign332(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign333(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign333(0 downto 0) <= BRAM_Dout_B(12 to 12);
  BRAM_Din_B(12 to 12) <= pgassign334(0 downto 0);
  pgassign335(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign335(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign335(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign335(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign336(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign336(0 downto 0) <= BRAM_Dout_A(13 to 13);
  BRAM_Din_A(13 to 13) <= pgassign337(0 downto 0);
  pgassign338(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign338(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign338(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign338(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign339(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign339(0 downto 0) <= BRAM_Dout_B(13 to 13);
  BRAM_Din_B(13 to 13) <= pgassign340(0 downto 0);
  pgassign341(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign341(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign341(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign341(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign342(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign342(0 downto 0) <= BRAM_Dout_A(14 to 14);
  BRAM_Din_A(14 to 14) <= pgassign343(0 downto 0);
  pgassign344(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign344(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign344(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign344(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign345(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign345(0 downto 0) <= BRAM_Dout_B(14 to 14);
  BRAM_Din_B(14 to 14) <= pgassign346(0 downto 0);
  pgassign347(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign347(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign347(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign347(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign348(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign348(0 downto 0) <= BRAM_Dout_A(15 to 15);
  BRAM_Din_A(15 to 15) <= pgassign349(0 downto 0);
  pgassign350(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign350(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign350(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign350(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign351(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign351(0 downto 0) <= BRAM_Dout_B(15 to 15);
  BRAM_Din_B(15 to 15) <= pgassign352(0 downto 0);
  pgassign353(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign353(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign353(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign353(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign354(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign354(0 downto 0) <= BRAM_Dout_A(16 to 16);
  BRAM_Din_A(16 to 16) <= pgassign355(0 downto 0);
  pgassign356(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign356(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign356(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign356(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign357(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign357(0 downto 0) <= BRAM_Dout_B(16 to 16);
  BRAM_Din_B(16 to 16) <= pgassign358(0 downto 0);
  pgassign359(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign359(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign359(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign359(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign360(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign360(0 downto 0) <= BRAM_Dout_A(17 to 17);
  BRAM_Din_A(17 to 17) <= pgassign361(0 downto 0);
  pgassign362(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign362(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign362(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign362(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign363(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign363(0 downto 0) <= BRAM_Dout_B(17 to 17);
  BRAM_Din_B(17 to 17) <= pgassign364(0 downto 0);
  pgassign365(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign365(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign365(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign365(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign366(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign366(0 downto 0) <= BRAM_Dout_A(18 to 18);
  BRAM_Din_A(18 to 18) <= pgassign367(0 downto 0);
  pgassign368(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign368(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign368(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign368(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign369(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign369(0 downto 0) <= BRAM_Dout_B(18 to 18);
  BRAM_Din_B(18 to 18) <= pgassign370(0 downto 0);
  pgassign371(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign371(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign371(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign371(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign372(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign372(0 downto 0) <= BRAM_Dout_A(19 to 19);
  BRAM_Din_A(19 to 19) <= pgassign373(0 downto 0);
  pgassign374(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign374(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign374(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign374(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign375(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign375(0 downto 0) <= BRAM_Dout_B(19 to 19);
  BRAM_Din_B(19 to 19) <= pgassign376(0 downto 0);
  pgassign377(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign377(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign377(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign377(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign378(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign378(0 downto 0) <= BRAM_Dout_A(20 to 20);
  BRAM_Din_A(20 to 20) <= pgassign379(0 downto 0);
  pgassign380(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign380(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign380(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign380(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign381(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign381(0 downto 0) <= BRAM_Dout_B(20 to 20);
  BRAM_Din_B(20 to 20) <= pgassign382(0 downto 0);
  pgassign383(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign383(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign383(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign383(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign384(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign384(0 downto 0) <= BRAM_Dout_A(21 to 21);
  BRAM_Din_A(21 to 21) <= pgassign385(0 downto 0);
  pgassign386(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign386(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign386(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign386(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign387(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign387(0 downto 0) <= BRAM_Dout_B(21 to 21);
  BRAM_Din_B(21 to 21) <= pgassign388(0 downto 0);
  pgassign389(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign389(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign389(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign389(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign390(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign390(0 downto 0) <= BRAM_Dout_A(22 to 22);
  BRAM_Din_A(22 to 22) <= pgassign391(0 downto 0);
  pgassign392(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign392(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign392(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign392(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign393(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign393(0 downto 0) <= BRAM_Dout_B(22 to 22);
  BRAM_Din_B(22 to 22) <= pgassign394(0 downto 0);
  pgassign395(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign395(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign395(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign395(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign396(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign396(0 downto 0) <= BRAM_Dout_A(23 to 23);
  BRAM_Din_A(23 to 23) <= pgassign397(0 downto 0);
  pgassign398(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign398(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign398(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign398(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign399(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign399(0 downto 0) <= BRAM_Dout_B(23 to 23);
  BRAM_Din_B(23 to 23) <= pgassign400(0 downto 0);
  pgassign401(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign401(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign401(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign401(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign402(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign402(0 downto 0) <= BRAM_Dout_A(24 to 24);
  BRAM_Din_A(24 to 24) <= pgassign403(0 downto 0);
  pgassign404(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign404(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign404(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign404(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign405(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign405(0 downto 0) <= BRAM_Dout_B(24 to 24);
  BRAM_Din_B(24 to 24) <= pgassign406(0 downto 0);
  pgassign407(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign407(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign407(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign407(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign408(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign408(0 downto 0) <= BRAM_Dout_A(25 to 25);
  BRAM_Din_A(25 to 25) <= pgassign409(0 downto 0);
  pgassign410(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign410(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign410(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign410(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign411(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign411(0 downto 0) <= BRAM_Dout_B(25 to 25);
  BRAM_Din_B(25 to 25) <= pgassign412(0 downto 0);
  pgassign413(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign413(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign413(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign413(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign414(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign414(0 downto 0) <= BRAM_Dout_A(26 to 26);
  BRAM_Din_A(26 to 26) <= pgassign415(0 downto 0);
  pgassign416(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign416(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign416(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign416(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign417(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign417(0 downto 0) <= BRAM_Dout_B(26 to 26);
  BRAM_Din_B(26 to 26) <= pgassign418(0 downto 0);
  pgassign419(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign419(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign419(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign419(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign420(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign420(0 downto 0) <= BRAM_Dout_A(27 to 27);
  BRAM_Din_A(27 to 27) <= pgassign421(0 downto 0);
  pgassign422(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign422(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign422(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign422(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign423(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign423(0 downto 0) <= BRAM_Dout_B(27 to 27);
  BRAM_Din_B(27 to 27) <= pgassign424(0 downto 0);
  pgassign425(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign425(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign425(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign425(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign426(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign426(0 downto 0) <= BRAM_Dout_A(28 to 28);
  BRAM_Din_A(28 to 28) <= pgassign427(0 downto 0);
  pgassign428(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign428(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign428(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign428(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign429(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign429(0 downto 0) <= BRAM_Dout_B(28 to 28);
  BRAM_Din_B(28 to 28) <= pgassign430(0 downto 0);
  pgassign431(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign431(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign431(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign431(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign432(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign432(0 downto 0) <= BRAM_Dout_A(29 to 29);
  BRAM_Din_A(29 to 29) <= pgassign433(0 downto 0);
  pgassign434(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign434(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign434(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign434(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign435(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign435(0 downto 0) <= BRAM_Dout_B(29 to 29);
  BRAM_Din_B(29 to 29) <= pgassign436(0 downto 0);
  pgassign437(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign437(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign437(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign437(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign438(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign438(0 downto 0) <= BRAM_Dout_A(30 to 30);
  BRAM_Din_A(30 to 30) <= pgassign439(0 downto 0);
  pgassign440(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign440(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign440(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign440(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign441(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign441(0 downto 0) <= BRAM_Dout_B(30 to 30);
  BRAM_Din_B(30 to 30) <= pgassign442(0 downto 0);
  pgassign443(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign443(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign443(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign443(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign444(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign444(0 downto 0) <= BRAM_Dout_A(31 to 31);
  BRAM_Din_A(31 to 31) <= pgassign445(0 downto 0);
  pgassign446(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign446(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign446(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign446(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign447(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign447(0 downto 0) <= BRAM_Dout_B(31 to 31);
  BRAM_Din_B(31 to 31) <= pgassign448(0 downto 0);
  pgassign449(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign449(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign449(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign449(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign450(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign450(0 downto 0) <= BRAM_Dout_A(32 to 32);
  BRAM_Din_A(32 to 32) <= pgassign451(0 downto 0);
  pgassign452(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign452(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign452(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign452(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign453(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign453(0 downto 0) <= BRAM_Dout_B(32 to 32);
  BRAM_Din_B(32 to 32) <= pgassign454(0 downto 0);
  pgassign455(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign455(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign455(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign455(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign456(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign456(0 downto 0) <= BRAM_Dout_A(33 to 33);
  BRAM_Din_A(33 to 33) <= pgassign457(0 downto 0);
  pgassign458(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign458(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign458(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign458(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign459(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign459(0 downto 0) <= BRAM_Dout_B(33 to 33);
  BRAM_Din_B(33 to 33) <= pgassign460(0 downto 0);
  pgassign461(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign461(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign461(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign461(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign462(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign462(0 downto 0) <= BRAM_Dout_A(34 to 34);
  BRAM_Din_A(34 to 34) <= pgassign463(0 downto 0);
  pgassign464(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign464(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign464(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign464(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign465(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign465(0 downto 0) <= BRAM_Dout_B(34 to 34);
  BRAM_Din_B(34 to 34) <= pgassign466(0 downto 0);
  pgassign467(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign467(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign467(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign467(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign468(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign468(0 downto 0) <= BRAM_Dout_A(35 to 35);
  BRAM_Din_A(35 to 35) <= pgassign469(0 downto 0);
  pgassign470(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign470(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign470(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign470(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign471(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign471(0 downto 0) <= BRAM_Dout_B(35 to 35);
  BRAM_Din_B(35 to 35) <= pgassign472(0 downto 0);
  pgassign473(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign473(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign473(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign473(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign474(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign474(0 downto 0) <= BRAM_Dout_A(36 to 36);
  BRAM_Din_A(36 to 36) <= pgassign475(0 downto 0);
  pgassign476(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign476(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign476(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign476(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign477(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign477(0 downto 0) <= BRAM_Dout_B(36 to 36);
  BRAM_Din_B(36 to 36) <= pgassign478(0 downto 0);
  pgassign479(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign479(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign479(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign479(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign480(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign480(0 downto 0) <= BRAM_Dout_A(37 to 37);
  BRAM_Din_A(37 to 37) <= pgassign481(0 downto 0);
  pgassign482(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign482(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign482(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign482(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign483(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign483(0 downto 0) <= BRAM_Dout_B(37 to 37);
  BRAM_Din_B(37 to 37) <= pgassign484(0 downto 0);
  pgassign485(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign485(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign485(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign485(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign486(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign486(0 downto 0) <= BRAM_Dout_A(38 to 38);
  BRAM_Din_A(38 to 38) <= pgassign487(0 downto 0);
  pgassign488(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign488(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign488(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign488(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign489(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign489(0 downto 0) <= BRAM_Dout_B(38 to 38);
  BRAM_Din_B(38 to 38) <= pgassign490(0 downto 0);
  pgassign491(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign491(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign491(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign491(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign492(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign492(0 downto 0) <= BRAM_Dout_A(39 to 39);
  BRAM_Din_A(39 to 39) <= pgassign493(0 downto 0);
  pgassign494(3 downto 3) <= BRAM_WEN_A(4 to 4);
  pgassign494(2 downto 2) <= BRAM_WEN_A(4 to 4);
  pgassign494(1 downto 1) <= BRAM_WEN_A(4 to 4);
  pgassign494(0 downto 0) <= BRAM_WEN_A(4 to 4);
  pgassign495(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign495(0 downto 0) <= BRAM_Dout_B(39 to 39);
  BRAM_Din_B(39 to 39) <= pgassign496(0 downto 0);
  pgassign497(3 downto 3) <= BRAM_WEN_B(4 to 4);
  pgassign497(2 downto 2) <= BRAM_WEN_B(4 to 4);
  pgassign497(1 downto 1) <= BRAM_WEN_B(4 to 4);
  pgassign497(0 downto 0) <= BRAM_WEN_B(4 to 4);
  pgassign498(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign498(0 downto 0) <= BRAM_Dout_A(40 to 40);
  BRAM_Din_A(40 to 40) <= pgassign499(0 downto 0);
  pgassign500(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign500(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign500(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign500(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign501(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign501(0 downto 0) <= BRAM_Dout_B(40 to 40);
  BRAM_Din_B(40 to 40) <= pgassign502(0 downto 0);
  pgassign503(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign503(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign503(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign503(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign504(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign504(0 downto 0) <= BRAM_Dout_A(41 to 41);
  BRAM_Din_A(41 to 41) <= pgassign505(0 downto 0);
  pgassign506(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign506(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign506(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign506(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign507(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign507(0 downto 0) <= BRAM_Dout_B(41 to 41);
  BRAM_Din_B(41 to 41) <= pgassign508(0 downto 0);
  pgassign509(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign509(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign509(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign509(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign510(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign510(0 downto 0) <= BRAM_Dout_A(42 to 42);
  BRAM_Din_A(42 to 42) <= pgassign511(0 downto 0);
  pgassign512(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign512(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign512(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign512(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign513(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign513(0 downto 0) <= BRAM_Dout_B(42 to 42);
  BRAM_Din_B(42 to 42) <= pgassign514(0 downto 0);
  pgassign515(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign515(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign515(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign515(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign516(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign516(0 downto 0) <= BRAM_Dout_A(43 to 43);
  BRAM_Din_A(43 to 43) <= pgassign517(0 downto 0);
  pgassign518(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign518(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign518(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign518(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign519(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign519(0 downto 0) <= BRAM_Dout_B(43 to 43);
  BRAM_Din_B(43 to 43) <= pgassign520(0 downto 0);
  pgassign521(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign521(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign521(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign521(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign522(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign522(0 downto 0) <= BRAM_Dout_A(44 to 44);
  BRAM_Din_A(44 to 44) <= pgassign523(0 downto 0);
  pgassign524(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign524(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign524(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign524(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign525(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign525(0 downto 0) <= BRAM_Dout_B(44 to 44);
  BRAM_Din_B(44 to 44) <= pgassign526(0 downto 0);
  pgassign527(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign527(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign527(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign527(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign528(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign528(0 downto 0) <= BRAM_Dout_A(45 to 45);
  BRAM_Din_A(45 to 45) <= pgassign529(0 downto 0);
  pgassign530(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign530(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign530(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign530(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign531(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign531(0 downto 0) <= BRAM_Dout_B(45 to 45);
  BRAM_Din_B(45 to 45) <= pgassign532(0 downto 0);
  pgassign533(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign533(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign533(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign533(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign534(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign534(0 downto 0) <= BRAM_Dout_A(46 to 46);
  BRAM_Din_A(46 to 46) <= pgassign535(0 downto 0);
  pgassign536(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign536(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign536(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign536(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign537(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign537(0 downto 0) <= BRAM_Dout_B(46 to 46);
  BRAM_Din_B(46 to 46) <= pgassign538(0 downto 0);
  pgassign539(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign539(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign539(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign539(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign540(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign540(0 downto 0) <= BRAM_Dout_A(47 to 47);
  BRAM_Din_A(47 to 47) <= pgassign541(0 downto 0);
  pgassign542(3 downto 3) <= BRAM_WEN_A(5 to 5);
  pgassign542(2 downto 2) <= BRAM_WEN_A(5 to 5);
  pgassign542(1 downto 1) <= BRAM_WEN_A(5 to 5);
  pgassign542(0 downto 0) <= BRAM_WEN_A(5 to 5);
  pgassign543(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign543(0 downto 0) <= BRAM_Dout_B(47 to 47);
  BRAM_Din_B(47 to 47) <= pgassign544(0 downto 0);
  pgassign545(3 downto 3) <= BRAM_WEN_B(5 to 5);
  pgassign545(2 downto 2) <= BRAM_WEN_B(5 to 5);
  pgassign545(1 downto 1) <= BRAM_WEN_B(5 to 5);
  pgassign545(0 downto 0) <= BRAM_WEN_B(5 to 5);
  pgassign546(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign546(0 downto 0) <= BRAM_Dout_A(48 to 48);
  BRAM_Din_A(48 to 48) <= pgassign547(0 downto 0);
  pgassign548(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign548(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign548(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign548(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign549(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign549(0 downto 0) <= BRAM_Dout_B(48 to 48);
  BRAM_Din_B(48 to 48) <= pgassign550(0 downto 0);
  pgassign551(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign551(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign551(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign551(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign552(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign552(0 downto 0) <= BRAM_Dout_A(49 to 49);
  BRAM_Din_A(49 to 49) <= pgassign553(0 downto 0);
  pgassign554(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign554(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign554(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign554(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign555(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign555(0 downto 0) <= BRAM_Dout_B(49 to 49);
  BRAM_Din_B(49 to 49) <= pgassign556(0 downto 0);
  pgassign557(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign557(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign557(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign557(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign558(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign558(0 downto 0) <= BRAM_Dout_A(50 to 50);
  BRAM_Din_A(50 to 50) <= pgassign559(0 downto 0);
  pgassign560(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign560(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign560(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign560(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign561(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign561(0 downto 0) <= BRAM_Dout_B(50 to 50);
  BRAM_Din_B(50 to 50) <= pgassign562(0 downto 0);
  pgassign563(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign563(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign563(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign563(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign564(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign564(0 downto 0) <= BRAM_Dout_A(51 to 51);
  BRAM_Din_A(51 to 51) <= pgassign565(0 downto 0);
  pgassign566(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign566(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign566(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign566(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign567(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign567(0 downto 0) <= BRAM_Dout_B(51 to 51);
  BRAM_Din_B(51 to 51) <= pgassign568(0 downto 0);
  pgassign569(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign569(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign569(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign569(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign570(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign570(0 downto 0) <= BRAM_Dout_A(52 to 52);
  BRAM_Din_A(52 to 52) <= pgassign571(0 downto 0);
  pgassign572(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign572(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign572(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign572(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign573(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign573(0 downto 0) <= BRAM_Dout_B(52 to 52);
  BRAM_Din_B(52 to 52) <= pgassign574(0 downto 0);
  pgassign575(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign575(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign575(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign575(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign576(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign576(0 downto 0) <= BRAM_Dout_A(53 to 53);
  BRAM_Din_A(53 to 53) <= pgassign577(0 downto 0);
  pgassign578(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign578(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign578(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign578(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign579(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign579(0 downto 0) <= BRAM_Dout_B(53 to 53);
  BRAM_Din_B(53 to 53) <= pgassign580(0 downto 0);
  pgassign581(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign581(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign581(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign581(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign582(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign582(0 downto 0) <= BRAM_Dout_A(54 to 54);
  BRAM_Din_A(54 to 54) <= pgassign583(0 downto 0);
  pgassign584(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign584(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign584(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign584(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign585(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign585(0 downto 0) <= BRAM_Dout_B(54 to 54);
  BRAM_Din_B(54 to 54) <= pgassign586(0 downto 0);
  pgassign587(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign587(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign587(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign587(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign588(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign588(0 downto 0) <= BRAM_Dout_A(55 to 55);
  BRAM_Din_A(55 to 55) <= pgassign589(0 downto 0);
  pgassign590(3 downto 3) <= BRAM_WEN_A(6 to 6);
  pgassign590(2 downto 2) <= BRAM_WEN_A(6 to 6);
  pgassign590(1 downto 1) <= BRAM_WEN_A(6 to 6);
  pgassign590(0 downto 0) <= BRAM_WEN_A(6 to 6);
  pgassign591(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign591(0 downto 0) <= BRAM_Dout_B(55 to 55);
  BRAM_Din_B(55 to 55) <= pgassign592(0 downto 0);
  pgassign593(3 downto 3) <= BRAM_WEN_B(6 to 6);
  pgassign593(2 downto 2) <= BRAM_WEN_B(6 to 6);
  pgassign593(1 downto 1) <= BRAM_WEN_B(6 to 6);
  pgassign593(0 downto 0) <= BRAM_WEN_B(6 to 6);
  pgassign594(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign594(0 downto 0) <= BRAM_Dout_A(56 to 56);
  BRAM_Din_A(56 to 56) <= pgassign595(0 downto 0);
  pgassign596(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign596(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign596(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign596(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign597(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign597(0 downto 0) <= BRAM_Dout_B(56 to 56);
  BRAM_Din_B(56 to 56) <= pgassign598(0 downto 0);
  pgassign599(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign599(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign599(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign599(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign600(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign600(0 downto 0) <= BRAM_Dout_A(57 to 57);
  BRAM_Din_A(57 to 57) <= pgassign601(0 downto 0);
  pgassign602(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign602(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign602(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign602(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign603(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign603(0 downto 0) <= BRAM_Dout_B(57 to 57);
  BRAM_Din_B(57 to 57) <= pgassign604(0 downto 0);
  pgassign605(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign605(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign605(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign605(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign606(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign606(0 downto 0) <= BRAM_Dout_A(58 to 58);
  BRAM_Din_A(58 to 58) <= pgassign607(0 downto 0);
  pgassign608(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign608(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign608(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign608(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign609(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign609(0 downto 0) <= BRAM_Dout_B(58 to 58);
  BRAM_Din_B(58 to 58) <= pgassign610(0 downto 0);
  pgassign611(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign611(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign611(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign611(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign612(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign612(0 downto 0) <= BRAM_Dout_A(59 to 59);
  BRAM_Din_A(59 to 59) <= pgassign613(0 downto 0);
  pgassign614(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign614(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign614(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign614(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign615(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign615(0 downto 0) <= BRAM_Dout_B(59 to 59);
  BRAM_Din_B(59 to 59) <= pgassign616(0 downto 0);
  pgassign617(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign617(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign617(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign617(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign618(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign618(0 downto 0) <= BRAM_Dout_A(60 to 60);
  BRAM_Din_A(60 to 60) <= pgassign619(0 downto 0);
  pgassign620(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign620(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign620(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign620(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign621(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign621(0 downto 0) <= BRAM_Dout_B(60 to 60);
  BRAM_Din_B(60 to 60) <= pgassign622(0 downto 0);
  pgassign623(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign623(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign623(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign623(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign624(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign624(0 downto 0) <= BRAM_Dout_A(61 to 61);
  BRAM_Din_A(61 to 61) <= pgassign625(0 downto 0);
  pgassign626(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign626(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign626(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign626(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign627(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign627(0 downto 0) <= BRAM_Dout_B(61 to 61);
  BRAM_Din_B(61 to 61) <= pgassign628(0 downto 0);
  pgassign629(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign629(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign629(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign629(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign630(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign630(0 downto 0) <= BRAM_Dout_A(62 to 62);
  BRAM_Din_A(62 to 62) <= pgassign631(0 downto 0);
  pgassign632(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign632(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign632(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign632(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign633(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign633(0 downto 0) <= BRAM_Dout_B(62 to 62);
  BRAM_Din_B(62 to 62) <= pgassign634(0 downto 0);
  pgassign635(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign635(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign635(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign635(0 downto 0) <= BRAM_WEN_B(7 to 7);
  pgassign636(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign636(0 downto 0) <= BRAM_Dout_A(63 to 63);
  BRAM_Din_A(63 to 63) <= pgassign637(0 downto 0);
  pgassign638(3 downto 3) <= BRAM_WEN_A(7 to 7);
  pgassign638(2 downto 2) <= BRAM_WEN_A(7 to 7);
  pgassign638(1 downto 1) <= BRAM_WEN_A(7 to 7);
  pgassign638(0 downto 0) <= BRAM_WEN_A(7 to 7);
  pgassign639(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign639(0 downto 0) <= BRAM_Dout_B(63 to 63);
  BRAM_Din_B(63 to 63) <= pgassign640(0 downto 0);
  pgassign641(3 downto 3) <= BRAM_WEN_B(7 to 7);
  pgassign641(2 downto 2) <= BRAM_WEN_B(7 to 7);
  pgassign641(1 downto 1) <= BRAM_WEN_B(7 to 7);
  pgassign641(0 downto 0) <= BRAM_WEN_B(7 to 7);
  net_gnd0 <= '0';
  net_gnd4(3 downto 0) <= B"0000";

  ramb16_0 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_0.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_0,
      CLKA => BRAM_Clk_A,
      DIA => pgassign2,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign3,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_0,
      CLKB => BRAM_Clk_B,
      DIB => pgassign4,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign5
    );

  ramb16_1 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_1.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_1,
      CLKA => BRAM_Clk_A,
      DIA => pgassign6,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign7,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_1,
      CLKB => BRAM_Clk_B,
      DIB => pgassign8,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign9
    );

  ramb16_2 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_2.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_2,
      CLKA => BRAM_Clk_A,
      DIA => pgassign10,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign11,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_2,
      CLKB => BRAM_Clk_B,
      DIB => pgassign12,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign13
    );

  ramb16_3 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_3.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_3,
      CLKA => BRAM_Clk_A,
      DIA => pgassign14,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign15,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_3,
      CLKB => BRAM_Clk_B,
      DIB => pgassign16,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign17
    );

  ramb16_4 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_4.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_4,
      CLKA => BRAM_Clk_A,
      DIA => pgassign18,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign19,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_4,
      CLKB => BRAM_Clk_B,
      DIB => pgassign20,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign21
    );

  ramb16_5 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_5.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_5,
      CLKA => BRAM_Clk_A,
      DIA => pgassign22,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign23,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_5,
      CLKB => BRAM_Clk_B,
      DIB => pgassign24,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign25
    );

  ramb16_6 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_6.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_6,
      CLKA => BRAM_Clk_A,
      DIA => pgassign26,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign27,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_6,
      CLKB => BRAM_Clk_B,
      DIB => pgassign28,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign29
    );

  ramb16_7 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_7.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_7,
      CLKA => BRAM_Clk_A,
      DIA => pgassign30,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign31,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_7,
      CLKB => BRAM_Clk_B,
      DIB => pgassign32,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign33
    );

  ramb16_8 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_8.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_8,
      CLKA => BRAM_Clk_A,
      DIA => pgassign34,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign35,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_8,
      CLKB => BRAM_Clk_B,
      DIB => pgassign36,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign37
    );

  ramb16_9 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_9.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_9,
      CLKA => BRAM_Clk_A,
      DIA => pgassign38,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign39,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_9,
      CLKB => BRAM_Clk_B,
      DIB => pgassign40,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign41
    );

  ramb16_10 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_10.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_10,
      CLKA => BRAM_Clk_A,
      DIA => pgassign42,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign43,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_10,
      CLKB => BRAM_Clk_B,
      DIB => pgassign44,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign45
    );

  ramb16_11 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_11.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_11,
      CLKA => BRAM_Clk_A,
      DIA => pgassign46,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign47,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_11,
      CLKB => BRAM_Clk_B,
      DIB => pgassign48,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign49
    );

  ramb16_12 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_12.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_12,
      CLKA => BRAM_Clk_A,
      DIA => pgassign50,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign51,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_12,
      CLKB => BRAM_Clk_B,
      DIB => pgassign52,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign53
    );

  ramb16_13 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_13.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_13,
      CLKA => BRAM_Clk_A,
      DIA => pgassign54,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign55,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_13,
      CLKB => BRAM_Clk_B,
      DIB => pgassign56,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign57
    );

  ramb16_14 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_14.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_14,
      CLKA => BRAM_Clk_A,
      DIA => pgassign58,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign59,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_14,
      CLKB => BRAM_Clk_B,
      DIB => pgassign60,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign61
    );

  ramb16_15 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_15.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_15,
      CLKA => BRAM_Clk_A,
      DIA => pgassign62,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign63,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_15,
      CLKB => BRAM_Clk_B,
      DIB => pgassign64,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign65
    );

  ramb16_16 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_16.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_16,
      CLKA => BRAM_Clk_A,
      DIA => pgassign66,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign67,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_16,
      CLKB => BRAM_Clk_B,
      DIB => pgassign68,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign69
    );

  ramb16_17 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_17.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_17,
      CLKA => BRAM_Clk_A,
      DIA => pgassign70,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign71,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_17,
      CLKB => BRAM_Clk_B,
      DIB => pgassign72,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign73
    );

  ramb16_18 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_18.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_18,
      CLKA => BRAM_Clk_A,
      DIA => pgassign74,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign75,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_18,
      CLKB => BRAM_Clk_B,
      DIB => pgassign76,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign77
    );

  ramb16_19 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_19.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_19,
      CLKA => BRAM_Clk_A,
      DIA => pgassign78,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign79,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_19,
      CLKB => BRAM_Clk_B,
      DIB => pgassign80,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign81
    );

  ramb16_20 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_20.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_20,
      CLKA => BRAM_Clk_A,
      DIA => pgassign82,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign83,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_20,
      CLKB => BRAM_Clk_B,
      DIB => pgassign84,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign85
    );

  ramb16_21 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_21.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_21,
      CLKA => BRAM_Clk_A,
      DIA => pgassign86,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign87,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_21,
      CLKB => BRAM_Clk_B,
      DIB => pgassign88,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign89
    );

  ramb16_22 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_22.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_22,
      CLKA => BRAM_Clk_A,
      DIA => pgassign90,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign91,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_22,
      CLKB => BRAM_Clk_B,
      DIB => pgassign92,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign93
    );

  ramb16_23 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_23.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_23,
      CLKA => BRAM_Clk_A,
      DIA => pgassign94,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign95,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_23,
      CLKB => BRAM_Clk_B,
      DIB => pgassign96,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign97
    );

  ramb16_24 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_24.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_24,
      CLKA => BRAM_Clk_A,
      DIA => pgassign98,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign99,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_24,
      CLKB => BRAM_Clk_B,
      DIB => pgassign100,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign101
    );

  ramb16_25 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_25.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_25,
      CLKA => BRAM_Clk_A,
      DIA => pgassign102,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign103,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_25,
      CLKB => BRAM_Clk_B,
      DIB => pgassign104,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign105
    );

  ramb16_26 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_26.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_26,
      CLKA => BRAM_Clk_A,
      DIA => pgassign106,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign107,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_26,
      CLKB => BRAM_Clk_B,
      DIB => pgassign108,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign109
    );

  ramb16_27 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_27.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_27,
      CLKA => BRAM_Clk_A,
      DIA => pgassign110,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign111,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_27,
      CLKB => BRAM_Clk_B,
      DIB => pgassign112,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign113
    );

  ramb16_28 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_28.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_28,
      CLKA => BRAM_Clk_A,
      DIA => pgassign114,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign115,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_28,
      CLKB => BRAM_Clk_B,
      DIB => pgassign116,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign117
    );

  ramb16_29 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_29.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_29,
      CLKA => BRAM_Clk_A,
      DIA => pgassign118,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign119,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_29,
      CLKB => BRAM_Clk_B,
      DIB => pgassign120,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign121
    );

  ramb16_30 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_30.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_30,
      CLKA => BRAM_Clk_A,
      DIA => pgassign122,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign123,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_30,
      CLKB => BRAM_Clk_B,
      DIB => pgassign124,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign125
    );

  ramb16_31 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_31.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_31,
      CLKA => BRAM_Clk_A,
      DIA => pgassign126,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign127,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_31,
      CLKB => BRAM_Clk_B,
      DIB => pgassign128,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign129
    );

  ramb16_32 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_32.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_32,
      CLKA => BRAM_Clk_A,
      DIA => pgassign130,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign131,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_32,
      CLKB => BRAM_Clk_B,
      DIB => pgassign132,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign133
    );

  ramb16_33 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_33.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_33,
      CLKA => BRAM_Clk_A,
      DIA => pgassign134,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign135,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_33,
      CLKB => BRAM_Clk_B,
      DIB => pgassign136,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign137
    );

  ramb16_34 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_34.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_34,
      CLKA => BRAM_Clk_A,
      DIA => pgassign138,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign139,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_34,
      CLKB => BRAM_Clk_B,
      DIB => pgassign140,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign141
    );

  ramb16_35 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_35.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_35,
      CLKA => BRAM_Clk_A,
      DIA => pgassign142,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign143,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_35,
      CLKB => BRAM_Clk_B,
      DIB => pgassign144,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign145
    );

  ramb16_36 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_36.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_36,
      CLKA => BRAM_Clk_A,
      DIA => pgassign146,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign147,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_36,
      CLKB => BRAM_Clk_B,
      DIB => pgassign148,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign149
    );

  ramb16_37 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_37.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_37,
      CLKA => BRAM_Clk_A,
      DIA => pgassign150,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign151,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_37,
      CLKB => BRAM_Clk_B,
      DIB => pgassign152,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign153
    );

  ramb16_38 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_38.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_38,
      CLKA => BRAM_Clk_A,
      DIA => pgassign154,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign155,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_38,
      CLKB => BRAM_Clk_B,
      DIB => pgassign156,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign157
    );

  ramb16_39 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_39.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_39,
      CLKA => BRAM_Clk_A,
      DIA => pgassign158,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign159,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_39,
      CLKB => BRAM_Clk_B,
      DIB => pgassign160,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign161
    );

  ramb16_40 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_40.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_40,
      CLKA => BRAM_Clk_A,
      DIA => pgassign162,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign163,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_40,
      CLKB => BRAM_Clk_B,
      DIB => pgassign164,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign165
    );

  ramb16_41 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_41.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_41,
      CLKA => BRAM_Clk_A,
      DIA => pgassign166,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign167,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_41,
      CLKB => BRAM_Clk_B,
      DIB => pgassign168,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign169
    );

  ramb16_42 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_42.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_42,
      CLKA => BRAM_Clk_A,
      DIA => pgassign170,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign171,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_42,
      CLKB => BRAM_Clk_B,
      DIB => pgassign172,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign173
    );

  ramb16_43 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_43.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_43,
      CLKA => BRAM_Clk_A,
      DIA => pgassign174,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign175,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_43,
      CLKB => BRAM_Clk_B,
      DIB => pgassign176,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign177
    );

  ramb16_44 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_44.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_44,
      CLKA => BRAM_Clk_A,
      DIA => pgassign178,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign179,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_44,
      CLKB => BRAM_Clk_B,
      DIB => pgassign180,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign181
    );

  ramb16_45 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_45.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_45,
      CLKA => BRAM_Clk_A,
      DIA => pgassign182,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign183,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_45,
      CLKB => BRAM_Clk_B,
      DIB => pgassign184,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign185
    );

  ramb16_46 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_46.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_46,
      CLKA => BRAM_Clk_A,
      DIA => pgassign186,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign187,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_46,
      CLKB => BRAM_Clk_B,
      DIB => pgassign188,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign189
    );

  ramb16_47 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_47.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_47,
      CLKA => BRAM_Clk_A,
      DIA => pgassign190,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign191,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_47,
      CLKB => BRAM_Clk_B,
      DIB => pgassign192,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign193
    );

  ramb16_48 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_48.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_48,
      CLKA => BRAM_Clk_A,
      DIA => pgassign194,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign195,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_48,
      CLKB => BRAM_Clk_B,
      DIB => pgassign196,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign197
    );

  ramb16_49 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_49.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_49,
      CLKA => BRAM_Clk_A,
      DIA => pgassign198,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign199,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_49,
      CLKB => BRAM_Clk_B,
      DIB => pgassign200,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign201
    );

  ramb16_50 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_50.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_50,
      CLKA => BRAM_Clk_A,
      DIA => pgassign202,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign203,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_50,
      CLKB => BRAM_Clk_B,
      DIB => pgassign204,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign205
    );

  ramb16_51 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_51.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_51,
      CLKA => BRAM_Clk_A,
      DIA => pgassign206,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign207,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_51,
      CLKB => BRAM_Clk_B,
      DIB => pgassign208,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign209
    );

  ramb16_52 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_52.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_52,
      CLKA => BRAM_Clk_A,
      DIA => pgassign210,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign211,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_52,
      CLKB => BRAM_Clk_B,
      DIB => pgassign212,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign213
    );

  ramb16_53 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_53.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_53,
      CLKA => BRAM_Clk_A,
      DIA => pgassign214,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign215,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_53,
      CLKB => BRAM_Clk_B,
      DIB => pgassign216,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign217
    );

  ramb16_54 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_54.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_54,
      CLKA => BRAM_Clk_A,
      DIA => pgassign218,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign219,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_54,
      CLKB => BRAM_Clk_B,
      DIB => pgassign220,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign221
    );

  ramb16_55 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_55.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_55,
      CLKA => BRAM_Clk_A,
      DIA => pgassign222,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign223,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_55,
      CLKB => BRAM_Clk_B,
      DIB => pgassign224,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign225
    );

  ramb16_56 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_56.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_56,
      CLKA => BRAM_Clk_A,
      DIA => pgassign226,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign227,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_56,
      CLKB => BRAM_Clk_B,
      DIB => pgassign228,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign229
    );

  ramb16_57 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_57.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_57,
      CLKA => BRAM_Clk_A,
      DIA => pgassign230,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign231,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_57,
      CLKB => BRAM_Clk_B,
      DIB => pgassign232,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign233
    );

  ramb16_58 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_58.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_58,
      CLKA => BRAM_Clk_A,
      DIA => pgassign234,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign235,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_58,
      CLKB => BRAM_Clk_B,
      DIB => pgassign236,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign237
    );

  ramb16_59 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_59.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_59,
      CLKA => BRAM_Clk_A,
      DIA => pgassign238,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign239,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_59,
      CLKB => BRAM_Clk_B,
      DIB => pgassign240,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign241
    );

  ramb16_60 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_60.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_60,
      CLKA => BRAM_Clk_A,
      DIA => pgassign242,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign243,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_60,
      CLKB => BRAM_Clk_B,
      DIB => pgassign244,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign245
    );

  ramb16_61 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_61.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_61,
      CLKA => BRAM_Clk_A,
      DIA => pgassign246,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign247,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_61,
      CLKB => BRAM_Clk_B,
      DIB => pgassign248,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign249
    );

  ramb16_62 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_62.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_62,
      CLKA => BRAM_Clk_A,
      DIA => pgassign250,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign251,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_62,
      CLKB => BRAM_Clk_B,
      DIB => pgassign252,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign253
    );

  ramb16_63 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_63.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "LOWER",
      RAM_EXTENSION_B => "LOWER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => net_gnd0,
      CASCADEOUTA => CASCADEA_63,
      CLKA => BRAM_Clk_A,
      DIA => pgassign254,
      DIPA => net_gnd4,
      DOA => open,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign255,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => net_gnd0,
      CASCADEOUTB => CASCADEB_63,
      CLKB => BRAM_Clk_B,
      DIB => pgassign256,
      DIPB => net_gnd4,
      DOB => open,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign257
    );

  ramb16_64 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_64.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_0,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign258,
      DIPA => net_gnd4,
      DOA => pgassign259,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign260,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_0,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign261,
      DIPB => net_gnd4,
      DOB => pgassign262,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign263
    );

  ramb16_65 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_65.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_1,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign264,
      DIPA => net_gnd4,
      DOA => pgassign265,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign266,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_1,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign267,
      DIPB => net_gnd4,
      DOB => pgassign268,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign269
    );

  ramb16_66 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_66.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_2,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign270,
      DIPA => net_gnd4,
      DOA => pgassign271,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign272,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_2,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign273,
      DIPB => net_gnd4,
      DOB => pgassign274,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign275
    );

  ramb16_67 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_67.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_3,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign276,
      DIPA => net_gnd4,
      DOA => pgassign277,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign278,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_3,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign279,
      DIPB => net_gnd4,
      DOB => pgassign280,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign281
    );

  ramb16_68 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_68.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_4,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign282,
      DIPA => net_gnd4,
      DOA => pgassign283,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign284,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_4,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign285,
      DIPB => net_gnd4,
      DOB => pgassign286,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign287
    );

  ramb16_69 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_69.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_5,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign288,
      DIPA => net_gnd4,
      DOA => pgassign289,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign290,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_5,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign291,
      DIPB => net_gnd4,
      DOB => pgassign292,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign293
    );

  ramb16_70 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_70.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_6,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign294,
      DIPA => net_gnd4,
      DOA => pgassign295,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign296,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_6,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign297,
      DIPB => net_gnd4,
      DOB => pgassign298,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign299
    );

  ramb16_71 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_71.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_7,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign300,
      DIPA => net_gnd4,
      DOA => pgassign301,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign302,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_7,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign303,
      DIPB => net_gnd4,
      DOB => pgassign304,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign305
    );

  ramb16_72 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_72.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_8,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign306,
      DIPA => net_gnd4,
      DOA => pgassign307,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign308,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_8,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign309,
      DIPB => net_gnd4,
      DOB => pgassign310,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign311
    );

  ramb16_73 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_73.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_9,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign312,
      DIPA => net_gnd4,
      DOA => pgassign313,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign314,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_9,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign315,
      DIPB => net_gnd4,
      DOB => pgassign316,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign317
    );

  ramb16_74 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_74.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_10,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign318,
      DIPA => net_gnd4,
      DOA => pgassign319,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign320,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_10,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign321,
      DIPB => net_gnd4,
      DOB => pgassign322,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign323
    );

  ramb16_75 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_75.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_11,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign324,
      DIPA => net_gnd4,
      DOA => pgassign325,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign326,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_11,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign327,
      DIPB => net_gnd4,
      DOB => pgassign328,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign329
    );

  ramb16_76 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_76.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_12,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign330,
      DIPA => net_gnd4,
      DOA => pgassign331,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign332,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_12,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign333,
      DIPB => net_gnd4,
      DOB => pgassign334,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign335
    );

  ramb16_77 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_77.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_13,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign336,
      DIPA => net_gnd4,
      DOA => pgassign337,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign338,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_13,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign339,
      DIPB => net_gnd4,
      DOB => pgassign340,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign341
    );

  ramb16_78 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_78.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_14,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign342,
      DIPA => net_gnd4,
      DOA => pgassign343,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign344,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_14,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign345,
      DIPB => net_gnd4,
      DOB => pgassign346,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign347
    );

  ramb16_79 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_79.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_15,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign348,
      DIPA => net_gnd4,
      DOA => pgassign349,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign350,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_15,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign351,
      DIPB => net_gnd4,
      DOB => pgassign352,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign353
    );

  ramb16_80 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_80.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_16,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign354,
      DIPA => net_gnd4,
      DOA => pgassign355,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign356,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_16,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign357,
      DIPB => net_gnd4,
      DOB => pgassign358,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign359
    );

  ramb16_81 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_81.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_17,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign360,
      DIPA => net_gnd4,
      DOA => pgassign361,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign362,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_17,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign363,
      DIPB => net_gnd4,
      DOB => pgassign364,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign365
    );

  ramb16_82 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_82.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_18,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign366,
      DIPA => net_gnd4,
      DOA => pgassign367,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign368,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_18,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign369,
      DIPB => net_gnd4,
      DOB => pgassign370,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign371
    );

  ramb16_83 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_83.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_19,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign372,
      DIPA => net_gnd4,
      DOA => pgassign373,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign374,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_19,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign375,
      DIPB => net_gnd4,
      DOB => pgassign376,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign377
    );

  ramb16_84 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_84.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_20,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign378,
      DIPA => net_gnd4,
      DOA => pgassign379,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign380,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_20,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign381,
      DIPB => net_gnd4,
      DOB => pgassign382,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign383
    );

  ramb16_85 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_85.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_21,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign384,
      DIPA => net_gnd4,
      DOA => pgassign385,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign386,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_21,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign387,
      DIPB => net_gnd4,
      DOB => pgassign388,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign389
    );

  ramb16_86 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_86.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_22,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign390,
      DIPA => net_gnd4,
      DOA => pgassign391,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign392,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_22,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign393,
      DIPB => net_gnd4,
      DOB => pgassign394,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign395
    );

  ramb16_87 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_87.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_23,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign396,
      DIPA => net_gnd4,
      DOA => pgassign397,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign398,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_23,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign399,
      DIPB => net_gnd4,
      DOB => pgassign400,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign401
    );

  ramb16_88 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_88.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_24,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign402,
      DIPA => net_gnd4,
      DOA => pgassign403,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign404,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_24,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign405,
      DIPB => net_gnd4,
      DOB => pgassign406,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign407
    );

  ramb16_89 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_89.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_25,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign408,
      DIPA => net_gnd4,
      DOA => pgassign409,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign410,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_25,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign411,
      DIPB => net_gnd4,
      DOB => pgassign412,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign413
    );

  ramb16_90 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_90.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_26,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign414,
      DIPA => net_gnd4,
      DOA => pgassign415,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign416,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_26,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign417,
      DIPB => net_gnd4,
      DOB => pgassign418,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign419
    );

  ramb16_91 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_91.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_27,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign420,
      DIPA => net_gnd4,
      DOA => pgassign421,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign422,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_27,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign423,
      DIPB => net_gnd4,
      DOB => pgassign424,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign425
    );

  ramb16_92 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_92.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_28,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign426,
      DIPA => net_gnd4,
      DOA => pgassign427,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign428,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_28,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign429,
      DIPB => net_gnd4,
      DOB => pgassign430,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign431
    );

  ramb16_93 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_93.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_29,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign432,
      DIPA => net_gnd4,
      DOA => pgassign433,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign434,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_29,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign435,
      DIPB => net_gnd4,
      DOB => pgassign436,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign437
    );

  ramb16_94 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_94.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_30,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign438,
      DIPA => net_gnd4,
      DOA => pgassign439,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign440,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_30,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign441,
      DIPB => net_gnd4,
      DOB => pgassign442,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign443
    );

  ramb16_95 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_95.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_31,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign444,
      DIPA => net_gnd4,
      DOA => pgassign445,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign446,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_31,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign447,
      DIPB => net_gnd4,
      DOB => pgassign448,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign449
    );

  ramb16_96 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_96.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_32,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign450,
      DIPA => net_gnd4,
      DOA => pgassign451,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign452,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_32,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign453,
      DIPB => net_gnd4,
      DOB => pgassign454,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign455
    );

  ramb16_97 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_97.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_33,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign456,
      DIPA => net_gnd4,
      DOA => pgassign457,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign458,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_33,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign459,
      DIPB => net_gnd4,
      DOB => pgassign460,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign461
    );

  ramb16_98 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_98.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_34,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign462,
      DIPA => net_gnd4,
      DOA => pgassign463,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign464,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_34,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign465,
      DIPB => net_gnd4,
      DOB => pgassign466,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign467
    );

  ramb16_99 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_99.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_35,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign468,
      DIPA => net_gnd4,
      DOA => pgassign469,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign470,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_35,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign471,
      DIPB => net_gnd4,
      DOB => pgassign472,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign473
    );

  ramb16_100 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_100.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_36,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign474,
      DIPA => net_gnd4,
      DOA => pgassign475,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign476,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_36,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign477,
      DIPB => net_gnd4,
      DOB => pgassign478,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign479
    );

  ramb16_101 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_101.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_37,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign480,
      DIPA => net_gnd4,
      DOA => pgassign481,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign482,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_37,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign483,
      DIPB => net_gnd4,
      DOB => pgassign484,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign485
    );

  ramb16_102 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_102.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_38,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign486,
      DIPA => net_gnd4,
      DOA => pgassign487,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign488,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_38,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign489,
      DIPB => net_gnd4,
      DOB => pgassign490,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign491
    );

  ramb16_103 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_103.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_39,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign492,
      DIPA => net_gnd4,
      DOA => pgassign493,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign494,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_39,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign495,
      DIPB => net_gnd4,
      DOB => pgassign496,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign497
    );

  ramb16_104 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_104.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_40,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign498,
      DIPA => net_gnd4,
      DOA => pgassign499,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign500,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_40,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign501,
      DIPB => net_gnd4,
      DOB => pgassign502,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign503
    );

  ramb16_105 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_105.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_41,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign504,
      DIPA => net_gnd4,
      DOA => pgassign505,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign506,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_41,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign507,
      DIPB => net_gnd4,
      DOB => pgassign508,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign509
    );

  ramb16_106 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_106.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_42,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign510,
      DIPA => net_gnd4,
      DOA => pgassign511,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign512,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_42,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign513,
      DIPB => net_gnd4,
      DOB => pgassign514,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign515
    );

  ramb16_107 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_107.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_43,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign516,
      DIPA => net_gnd4,
      DOA => pgassign517,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign518,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_43,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign519,
      DIPB => net_gnd4,
      DOB => pgassign520,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign521
    );

  ramb16_108 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_108.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_44,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign522,
      DIPA => net_gnd4,
      DOA => pgassign523,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign524,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_44,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign525,
      DIPB => net_gnd4,
      DOB => pgassign526,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign527
    );

  ramb16_109 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_109.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_45,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign528,
      DIPA => net_gnd4,
      DOA => pgassign529,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign530,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_45,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign531,
      DIPB => net_gnd4,
      DOB => pgassign532,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign533
    );

  ramb16_110 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_110.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_46,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign534,
      DIPA => net_gnd4,
      DOA => pgassign535,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign536,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_46,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign537,
      DIPB => net_gnd4,
      DOB => pgassign538,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign539
    );

  ramb16_111 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_111.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_47,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign540,
      DIPA => net_gnd4,
      DOA => pgassign541,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign542,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_47,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign543,
      DIPB => net_gnd4,
      DOB => pgassign544,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign545
    );

  ramb16_112 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_112.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_48,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign546,
      DIPA => net_gnd4,
      DOA => pgassign547,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign548,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_48,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign549,
      DIPB => net_gnd4,
      DOB => pgassign550,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign551
    );

  ramb16_113 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_113.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_49,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign552,
      DIPA => net_gnd4,
      DOA => pgassign553,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign554,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_49,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign555,
      DIPB => net_gnd4,
      DOB => pgassign556,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign557
    );

  ramb16_114 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_114.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_50,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign558,
      DIPA => net_gnd4,
      DOA => pgassign559,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign560,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_50,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign561,
      DIPB => net_gnd4,
      DOB => pgassign562,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign563
    );

  ramb16_115 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_115.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_51,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign564,
      DIPA => net_gnd4,
      DOA => pgassign565,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign566,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_51,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign567,
      DIPB => net_gnd4,
      DOB => pgassign568,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign569
    );

  ramb16_116 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_116.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_52,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign570,
      DIPA => net_gnd4,
      DOA => pgassign571,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign572,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_52,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign573,
      DIPB => net_gnd4,
      DOB => pgassign574,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign575
    );

  ramb16_117 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_117.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_53,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign576,
      DIPA => net_gnd4,
      DOA => pgassign577,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign578,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_53,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign579,
      DIPB => net_gnd4,
      DOB => pgassign580,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign581
    );

  ramb16_118 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_118.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_54,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign582,
      DIPA => net_gnd4,
      DOA => pgassign583,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign584,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_54,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign585,
      DIPB => net_gnd4,
      DOB => pgassign586,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign587
    );

  ramb16_119 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_119.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_55,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign588,
      DIPA => net_gnd4,
      DOA => pgassign589,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign590,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_55,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign591,
      DIPB => net_gnd4,
      DOB => pgassign592,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign593
    );

  ramb16_120 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_120.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_56,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign594,
      DIPA => net_gnd4,
      DOA => pgassign595,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign596,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_56,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign597,
      DIPB => net_gnd4,
      DOB => pgassign598,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign599
    );

  ramb16_121 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_121.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_57,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign600,
      DIPA => net_gnd4,
      DOA => pgassign601,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign602,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_57,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign603,
      DIPB => net_gnd4,
      DOB => pgassign604,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign605
    );

  ramb16_122 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_122.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_58,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign606,
      DIPA => net_gnd4,
      DOA => pgassign607,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign608,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_58,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign609,
      DIPB => net_gnd4,
      DOB => pgassign610,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign611
    );

  ramb16_123 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_123.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_59,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign612,
      DIPA => net_gnd4,
      DOA => pgassign613,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign614,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_59,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign615,
      DIPB => net_gnd4,
      DOB => pgassign616,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign617
    );

  ramb16_124 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_124.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_60,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign618,
      DIPA => net_gnd4,
      DOA => pgassign619,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign620,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_60,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign621,
      DIPB => net_gnd4,
      DOB => pgassign622,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign623
    );

  ramb16_125 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_125.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_61,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign624,
      DIPA => net_gnd4,
      DOA => pgassign625,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign626,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_61,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign627,
      DIPB => net_gnd4,
      DOB => pgassign628,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign629
    );

  ramb16_126 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_126.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_62,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign630,
      DIPA => net_gnd4,
      DOA => pgassign631,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign632,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_62,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign633,
      DIPB => net_gnd4,
      DOB => pgassign634,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign635
    );

  ramb16_127 : RAMB16
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "plb_bram_if_cntlr_0_bram_combined_127.mem",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "UPPER",
      RAM_EXTENSION_B => "UPPER"
    )
    port map (
      ADDRA => BRAM_Addr_A(14 to 28),
      CASCADEINA => CASCADEA_63,
      CASCADEOUTA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign636,
      DIPA => net_gnd4,
      DOA => pgassign637,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign638,
      ADDRB => BRAM_Addr_B(14 to 28),
      CASCADEINB => CASCADEB_63,
      CASCADEOUTB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign639,
      DIPB => net_gnd4,
      DOB => pgassign640,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign641
    );

end architecture STRUCTURE;

